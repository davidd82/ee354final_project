module tictactoeboard_rom
	(
		input wire clk,
		input wire [8:0] row,
		input wire [9:0] col,
		output reg [11:0] color_data
	);

	(* rom_style = "block" *)

	//signal declaration
	reg [8:0] row_reg;
	reg [9:0] col_reg;

	always @(posedge clk)
		begin
		row_reg <= row;
		col_reg <= col;
		end

	always @(*) begin
		if(({row_reg, col_reg}>=19'b0000000000000000000) && ({row_reg, col_reg}<19'b0000000000011110000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0000000000011110000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0000000000011110001)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0000000000011110010)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0000000000011110011)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0000000000011110100)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0000000000011110101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0000000000011110110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0000000000011110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0000000000011111000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0000000000011111001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0000000000011111010)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0000000000011111011)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=19'b0000000000011111100) && ({row_reg, col_reg}<19'b0000000000110000110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=19'b0000000000110000110) && ({row_reg, col_reg}<19'b0000000000110001000)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0000000000110001000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0000000000110001001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0000000000110001010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0000000000110001011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0000000000110001100)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0000000000110001101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0000000000110001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0000000000110001111)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0000000000110010000)) color_data = 12'b110111011101;

		if(({row_reg, col_reg}>=19'b0000000000110010001) && ({row_reg, col_reg}<19'b0000000010011101110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0000000010011101110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0000000010011101111)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0000000010011110000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0000000010011110001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=19'b0000000010011110010) && ({row_reg, col_reg}<19'b0000000010011110110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000000010011110110) && ({row_reg, col_reg}<19'b0000000010011111000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0000000010011111000) && ({row_reg, col_reg}<19'b0000000010011111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0000000010011111010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0000000010011111011)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0000000010011111100)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=19'b0000000010011111101) && ({row_reg, col_reg}<19'b0000000010110000100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0000000010110000100)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0000000010110000101)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0000000010110000110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=19'b0000000010110000111) && ({row_reg, col_reg}<19'b0000000010110001010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000000010110001010) && ({row_reg, col_reg}<19'b0000000010110001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0000000010110001100) && ({row_reg, col_reg}<19'b0000000010110010000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0000000010110010000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0000000010110010001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0000000010110010010)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0000000010110010011) && ({row_reg, col_reg}<19'b0000000100011101101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0000000100011101101)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0000000100011101110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0000000100011101111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0000000100011110000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000000100011110001) && ({row_reg, col_reg}<19'b0000000100011110111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000000100011110111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0000000100011111000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000000100011111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000000100011111010) && ({row_reg, col_reg}<19'b0000000100011111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000000100011111100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0000000100011111101)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0000000100011111110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=19'b0000000100011111111) && ({row_reg, col_reg}<19'b0000000100110000011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0000000100110000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0000000100110000100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=19'b0000000100110000101) && ({row_reg, col_reg}<19'b0000000100110000111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0000000100110000111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000000100110001000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0000000100110001001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0000000100110001010) && ({row_reg, col_reg}<19'b0000000100110001101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000000100110001101) && ({row_reg, col_reg}<19'b0000000100110001111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0000000100110001111) && ({row_reg, col_reg}<19'b0000000100110010010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0000000100110010010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0000000100110010011)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0000000100110010100)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0000000100110010101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0000000100110010110)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0000000100110010111) && ({row_reg, col_reg}<19'b0000000110011101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0000000110011101100)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0000000110011101101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=19'b0000000110011101110) && ({row_reg, col_reg}<19'b0000000110011110000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0000000110011110000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0000000110011110001) && ({row_reg, col_reg}<19'b0000000110011111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0000000110011111011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0000000110011111100) && ({row_reg, col_reg}<19'b0000000110011111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0000000110011111110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0000000110011111111)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=19'b0000000110100000000) && ({row_reg, col_reg}<19'b0000000110110000010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0000000110110000010)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0000000110110000011)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0000000110110000100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000000110110000101) && ({row_reg, col_reg}<19'b0000000110110000111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000000110110000111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000000110110001000) && ({row_reg, col_reg}<19'b0000000110110010010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000000110110010010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0000000110110010011)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0000000110110010100)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0000000110110010101)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0000000110110010110) && ({row_reg, col_reg}<19'b0000001000011101011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0000001000011101011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0000001000011101100)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0000001000011101101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0000001000011101110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000001000011101111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000001000011110000) && ({row_reg, col_reg}<19'b0000001000011111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0000001000011111010) && ({row_reg, col_reg}<19'b0000001000011111101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0000001000011111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000001000011111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0000001000011111111)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0000001000100000000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=19'b0000001000100000001) && ({row_reg, col_reg}<19'b0000001000110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0000001000110000001)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0000001000110000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0000001000110000011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0000001000110000100) && ({row_reg, col_reg}<19'b0000001000110000110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000001000110000110) && ({row_reg, col_reg}<19'b0000001000110001000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0000001000110001000) && ({row_reg, col_reg}<19'b0000001000110001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000001000110001110) && ({row_reg, col_reg}<19'b0000001000110010011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0000001000110010011) && ({row_reg, col_reg}<19'b0000001000110010101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0000001000110010101)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=19'b0000001000110010110) && ({row_reg, col_reg}<19'b0000001010011101010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0000001010011101010)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0000001010011101011)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=19'b0000001010011101100) && ({row_reg, col_reg}<19'b0000001010011101111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000001010011101111) && ({row_reg, col_reg}<19'b0000001010011110001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0000001010011110001) && ({row_reg, col_reg}<19'b0000001010011110100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000001010011110100) && ({row_reg, col_reg}<19'b0000001010011110110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0000001010011110110) && ({row_reg, col_reg}<19'b0000001010011111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000001010011111011) && ({row_reg, col_reg}<19'b0000001010011111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0000001010011111101) && ({row_reg, col_reg}<19'b0000001010100000000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0000001010100000000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0000001010100000001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=19'b0000001010100000010) && ({row_reg, col_reg}<19'b0000001010110000000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0000001010110000000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0000001010110000001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0000001010110000010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000001010110000011) && ({row_reg, col_reg}<19'b0000001010110000111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0000001010110000111) && ({row_reg, col_reg}<19'b0000001010110001010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000001010110001010) && ({row_reg, col_reg}<19'b0000001010110010000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000001010110010000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000001010110010001) && ({row_reg, col_reg}<19'b0000001010110010011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000001010110010011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0000001010110010100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000001010110010101)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0000001010110010110)) color_data = 12'b110111011101;

		if(({row_reg, col_reg}>=19'b0000001010110010111) && ({row_reg, col_reg}<19'b0000001100011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0000001100011101000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0000001100011101001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0000001100011101010)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0000001100011101011)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=19'b0000001100011101100) && ({row_reg, col_reg}<19'b0000001100011101111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000001100011101111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000001100011110000) && ({row_reg, col_reg}<19'b0000001100011110101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000001100011110101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000001100011110110) && ({row_reg, col_reg}<19'b0000001100011111000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000001100011111000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000001100011111001) && ({row_reg, col_reg}<19'b0000001100011111011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0000001100011111011) && ({row_reg, col_reg}<19'b0000001100011111101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000001100011111101) && ({row_reg, col_reg}<19'b0000001100011111111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000001100011111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0000001100100000000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0000001100100000001)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0000001100100000010) && ({row_reg, col_reg}<19'b0000001100101111111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0000001100101111111)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0000001100110000000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0000001100110000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000001100110000010) && ({row_reg, col_reg}<19'b0000001100110000101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000001100110000101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0000001100110000110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000001100110000111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000001100110001000) && ({row_reg, col_reg}<19'b0000001100110001010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0000001100110001010) && ({row_reg, col_reg}<19'b0000001100110001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000001100110001110) && ({row_reg, col_reg}<19'b0000001100110010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0000001100110010001) && ({row_reg, col_reg}<19'b0000001100110010011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000001100110010011) && ({row_reg, col_reg}<19'b0000001100110010101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000001100110010101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0000001100110010110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0000001100110010111)) color_data = 12'b110111011101;

		if(({row_reg, col_reg}>=19'b0000001100110011000) && ({row_reg, col_reg}<19'b0000001110011101001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0000001110011101001)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0000001110011101010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0000001110011101011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0000001110011101100) && ({row_reg, col_reg}<19'b0000001110011101111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000001110011101111) && ({row_reg, col_reg}<19'b0000001110011110111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000001110011110111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000001110011111000) && ({row_reg, col_reg}<19'b0000001110011111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0000001110011111010) && ({row_reg, col_reg}<19'b0000001110011111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000001110011111100) && ({row_reg, col_reg}<19'b0000001110011111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000001110011111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000001110011111111) && ({row_reg, col_reg}<19'b0000001110100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000001110100000001)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0000001110100000010)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=19'b0000001110100000011) && ({row_reg, col_reg}<19'b0000001110101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0000001110101111110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0000001110101111111)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0000001110110000000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0000001110110000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000001110110000010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000001110110000011) && ({row_reg, col_reg}<19'b0000001110110000101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000001110110000101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000001110110000110) && ({row_reg, col_reg}<19'b0000001110110001001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0000001110110001001) && ({row_reg, col_reg}<19'b0000001110110001011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000001110110001011) && ({row_reg, col_reg}<19'b0000001110110010000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000001110110010000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000001110110010001) && ({row_reg, col_reg}<19'b0000001110110010100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000001110110010100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0000001110110010101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000001110110010110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0000001110110010111)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=19'b0000001110110011000) && ({row_reg, col_reg}<19'b0000010000011101001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0000010000011101001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0000010000011101010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0000010000011101011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000010000011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0000010000011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000010000011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000010000011101111) && ({row_reg, col_reg}<19'b0000010000100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000010000100000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0000010000100000010)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0000010000100000011) && ({row_reg, col_reg}<19'b0000010000101111111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0000010000101111111)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=19'b0000010000110000000) && ({row_reg, col_reg}<19'b0000010000110000011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000010000110000011) && ({row_reg, col_reg}<19'b0000010000110010010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000010000110010010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000010000110010011) && ({row_reg, col_reg}<19'b0000010000110010110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000010000110010110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0000010000110010111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0000010000110011000)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0000010000110011001) && ({row_reg, col_reg}<19'b0000010010011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0000010010011101000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0000010010011101001)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0000010010011101010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0000010010011101011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000010010011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000010010011101101) && ({row_reg, col_reg}<19'b0000010010100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000010010100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0000010010100000010)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=19'b0000010010100000011) && ({row_reg, col_reg}<19'b0000010010101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0000010010101111110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0000010010101111111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=19'b0000010010110000000) && ({row_reg, col_reg}<19'b0000010010110010000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000010010110010000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0000010010110010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000010010110010010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000010010110010011) && ({row_reg, col_reg}<19'b0000010010110010111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000010010110010111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0000010010110011000)) color_data = 12'b110111011101;

		if(({row_reg, col_reg}>=19'b0000010010110011001) && ({row_reg, col_reg}<19'b0000010100011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0000010100011101000)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0000010100011101001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0000010100011101010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0000010100011101011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000010100011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000010100011101101) && ({row_reg, col_reg}<19'b0000010100011101111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000010100011101111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000010100011110000) && ({row_reg, col_reg}<19'b0000010100100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000010100100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0000010100100000010)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=19'b0000010100100000011) && ({row_reg, col_reg}<19'b0000010100101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0000010100101111110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0000010100101111111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=19'b0000010100110000000) && ({row_reg, col_reg}<19'b0000010100110010000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000010100110010000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0000010100110010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000010100110010010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0000010100110010011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0000010100110010100) && ({row_reg, col_reg}<19'b0000010100110010110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0000010100110010110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000010100110010111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0000010100110011000)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=19'b0000010100110011001) && ({row_reg, col_reg}<19'b0000010110011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0000010110011101000)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0000010110011101001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=19'b0000010110011101010) && ({row_reg, col_reg}<19'b0000010110011101101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000010110011101101) && ({row_reg, col_reg}<19'b0000010110011101111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000010110011101111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000010110011110000) && ({row_reg, col_reg}<19'b0000010110100000000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0000010110100000000) && ({row_reg, col_reg}<19'b0000010110100000010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0000010110100000010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0000010110100000011)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=19'b0000010110100000100) && ({row_reg, col_reg}<19'b0000010110101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0000010110101111110)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0000010110101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000010110110000000) && ({row_reg, col_reg}<19'b0000010110110010010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000010110110010010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0000010110110010011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0000010110110010100) && ({row_reg, col_reg}<19'b0000010110110010110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0000010110110010110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000010110110010111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0000010110110011000)) color_data = 12'b101110111011;

		if(({row_reg, col_reg}>=19'b0000010110110011001) && ({row_reg, col_reg}<19'b0000011000011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0000011000011101000)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0000011000011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0000011000011101010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000011000011101011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000011000011101100) && ({row_reg, col_reg}<19'b0000011000100000000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0000011000100000000) && ({row_reg, col_reg}<19'b0000011000100000010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0000011000100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0000011000100000011)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=19'b0000011000100000100) && ({row_reg, col_reg}<19'b0000011000101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0000011000101111110)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0000011000101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000011000110000000) && ({row_reg, col_reg}<19'b0000011000110010010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000011000110010010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000011000110010011) && ({row_reg, col_reg}<19'b0000011000110010101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0000011000110010101) && ({row_reg, col_reg}<19'b0000011000110011000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0000011000110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0000011000110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0000011000110011010) && ({row_reg, col_reg}<19'b0000011010011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0000011010011101000)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0000011010011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000011010011101010) && ({row_reg, col_reg}<19'b0000011010011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000011010011101101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000011010011101110) && ({row_reg, col_reg}<19'b0000011010100000010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000011010100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0000011010100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0000011010100000100) && ({row_reg, col_reg}<19'b0000011010101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0000011010101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0000011010101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000011010110000000) && ({row_reg, col_reg}<19'b0000011010110010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0000011010110010001) && ({row_reg, col_reg}<19'b0000011010110010011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000011010110010011) && ({row_reg, col_reg}<19'b0000011010110010111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000011010110010111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0000011010110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0000011010110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0000011010110011010) && ({row_reg, col_reg}<19'b0000011100011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0000011100011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0000011100011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000011100011101010) && ({row_reg, col_reg}<19'b0000011100011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0000011100011101100) && ({row_reg, col_reg}<19'b0000011100011101111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000011100011101111) && ({row_reg, col_reg}<19'b0000011100100000010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000011100100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0000011100100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0000011100100000100) && ({row_reg, col_reg}<19'b0000011100101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0000011100101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=19'b0000011100101111111) && ({row_reg, col_reg}<19'b0000011100110000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000011100110000001) && ({row_reg, col_reg}<19'b0000011100110010011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000011100110010011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000011100110010100) && ({row_reg, col_reg}<19'b0000011100110010110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000011100110010110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0000011100110010111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000011100110011000)) color_data = 12'b101010101010;

		if(({row_reg, col_reg}>=19'b0000011100110011001) && ({row_reg, col_reg}<19'b0000011110011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0000011110011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=19'b0000011110011101001) && ({row_reg, col_reg}<19'b0000011110011101011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0000011110011101011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000011110011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000011110011101101) && ({row_reg, col_reg}<19'b0000011110100000010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000011110100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0000011110100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0000011110100000100) && ({row_reg, col_reg}<19'b0000011110101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0000011110101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0000011110101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000011110110000000) && ({row_reg, col_reg}<19'b0000011110110000111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000011110110000111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000011110110001000) && ({row_reg, col_reg}<19'b0000011110110010000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000011110110010000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000011110110010001) && ({row_reg, col_reg}<19'b0000011110110010011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0000011110110010011) && ({row_reg, col_reg}<19'b0000011110110010101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0000011110110010101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000011110110010110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0000011110110010111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000011110110011000)) color_data = 12'b101010101010;

		if(({row_reg, col_reg}>=19'b0000011110110011001) && ({row_reg, col_reg}<19'b0000100000011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0000100000011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0000100000011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000100000011101010) && ({row_reg, col_reg}<19'b0000100000011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000100000011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0000100000011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000100000011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000100000011101111) && ({row_reg, col_reg}<19'b0000100000100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000100000100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0000100000100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0000100000100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0000100000100000100) && ({row_reg, col_reg}<19'b0000100000101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0000100000101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0000100000101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000100000110000000) && ({row_reg, col_reg}<19'b0000100000110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000100000110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0000100000110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0000100000110011010) && ({row_reg, col_reg}<19'b0000100010011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0000100010011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0000100010011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000100010011101010) && ({row_reg, col_reg}<19'b0000100010011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000100010011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0000100010011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000100010011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000100010011101111) && ({row_reg, col_reg}<19'b0000100010100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000100010100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0000100010100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0000100010100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0000100010100000100) && ({row_reg, col_reg}<19'b0000100010101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0000100010101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0000100010101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000100010110000000) && ({row_reg, col_reg}<19'b0000100010110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000100010110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0000100010110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0000100010110011010) && ({row_reg, col_reg}<19'b0000100100011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0000100100011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0000100100011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000100100011101010) && ({row_reg, col_reg}<19'b0000100100011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000100100011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0000100100011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000100100011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000100100011101111) && ({row_reg, col_reg}<19'b0000100100100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000100100100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0000100100100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0000100100100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0000100100100000100) && ({row_reg, col_reg}<19'b0000100100101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0000100100101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0000100100101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000100100110000000) && ({row_reg, col_reg}<19'b0000100100110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000100100110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0000100100110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0000100100110011010) && ({row_reg, col_reg}<19'b0000100110011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0000100110011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0000100110011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000100110011101010) && ({row_reg, col_reg}<19'b0000100110011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000100110011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0000100110011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000100110011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000100110011101111) && ({row_reg, col_reg}<19'b0000100110100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000100110100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0000100110100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0000100110100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0000100110100000100) && ({row_reg, col_reg}<19'b0000100110101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0000100110101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0000100110101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000100110110000000) && ({row_reg, col_reg}<19'b0000100110110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000100110110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0000100110110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0000100110110011010) && ({row_reg, col_reg}<19'b0000101000011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0000101000011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0000101000011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000101000011101010) && ({row_reg, col_reg}<19'b0000101000011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000101000011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0000101000011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000101000011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000101000011101111) && ({row_reg, col_reg}<19'b0000101000100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000101000100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0000101000100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0000101000100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0000101000100000100) && ({row_reg, col_reg}<19'b0000101000101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0000101000101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0000101000101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000101000110000000) && ({row_reg, col_reg}<19'b0000101000110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000101000110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0000101000110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0000101000110011010) && ({row_reg, col_reg}<19'b0000101010011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0000101010011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0000101010011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000101010011101010) && ({row_reg, col_reg}<19'b0000101010011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000101010011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0000101010011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000101010011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000101010011101111) && ({row_reg, col_reg}<19'b0000101010100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000101010100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0000101010100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0000101010100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0000101010100000100) && ({row_reg, col_reg}<19'b0000101010101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0000101010101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0000101010101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000101010110000000) && ({row_reg, col_reg}<19'b0000101010110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000101010110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0000101010110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0000101010110011010) && ({row_reg, col_reg}<19'b0000101100011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0000101100011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0000101100011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000101100011101010) && ({row_reg, col_reg}<19'b0000101100011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000101100011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0000101100011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000101100011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000101100011101111) && ({row_reg, col_reg}<19'b0000101100100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000101100100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0000101100100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0000101100100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0000101100100000100) && ({row_reg, col_reg}<19'b0000101100101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0000101100101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0000101100101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000101100110000000) && ({row_reg, col_reg}<19'b0000101100110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000101100110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0000101100110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0000101100110011010) && ({row_reg, col_reg}<19'b0000101110011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0000101110011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0000101110011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000101110011101010) && ({row_reg, col_reg}<19'b0000101110011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000101110011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0000101110011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000101110011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000101110011101111) && ({row_reg, col_reg}<19'b0000101110100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000101110100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0000101110100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0000101110100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0000101110100000100) && ({row_reg, col_reg}<19'b0000101110101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0000101110101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0000101110101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000101110110000000) && ({row_reg, col_reg}<19'b0000101110110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000101110110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0000101110110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0000101110110011010) && ({row_reg, col_reg}<19'b0000110000011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0000110000011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0000110000011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000110000011101010) && ({row_reg, col_reg}<19'b0000110000011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000110000011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0000110000011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000110000011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000110000011101111) && ({row_reg, col_reg}<19'b0000110000100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000110000100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0000110000100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0000110000100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0000110000100000100) && ({row_reg, col_reg}<19'b0000110000101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0000110000101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0000110000101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000110000110000000) && ({row_reg, col_reg}<19'b0000110000110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000110000110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0000110000110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0000110000110011010) && ({row_reg, col_reg}<19'b0000110010011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0000110010011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0000110010011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000110010011101010) && ({row_reg, col_reg}<19'b0000110010011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000110010011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0000110010011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000110010011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000110010011101111) && ({row_reg, col_reg}<19'b0000110010100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000110010100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0000110010100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0000110010100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0000110010100000100) && ({row_reg, col_reg}<19'b0000110010101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0000110010101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0000110010101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000110010110000000) && ({row_reg, col_reg}<19'b0000110010110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000110010110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0000110010110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0000110010110011010) && ({row_reg, col_reg}<19'b0000110100011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0000110100011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0000110100011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000110100011101010) && ({row_reg, col_reg}<19'b0000110100011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000110100011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0000110100011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000110100011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000110100011101111) && ({row_reg, col_reg}<19'b0000110100100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000110100100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0000110100100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0000110100100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0000110100100000100) && ({row_reg, col_reg}<19'b0000110100101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0000110100101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0000110100101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000110100110000000) && ({row_reg, col_reg}<19'b0000110100110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000110100110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0000110100110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0000110100110011010) && ({row_reg, col_reg}<19'b0000110110011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0000110110011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0000110110011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000110110011101010) && ({row_reg, col_reg}<19'b0000110110011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000110110011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0000110110011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000110110011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000110110011101111) && ({row_reg, col_reg}<19'b0000110110100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000110110100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0000110110100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0000110110100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0000110110100000100) && ({row_reg, col_reg}<19'b0000110110101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0000110110101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0000110110101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000110110110000000) && ({row_reg, col_reg}<19'b0000110110110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000110110110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0000110110110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0000110110110011010) && ({row_reg, col_reg}<19'b0000111000011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0000111000011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0000111000011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000111000011101010) && ({row_reg, col_reg}<19'b0000111000011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000111000011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0000111000011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000111000011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000111000011101111) && ({row_reg, col_reg}<19'b0000111000100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000111000100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0000111000100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0000111000100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0000111000100000100) && ({row_reg, col_reg}<19'b0000111000101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0000111000101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0000111000101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000111000110000000) && ({row_reg, col_reg}<19'b0000111000110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000111000110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0000111000110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0000111000110011010) && ({row_reg, col_reg}<19'b0000111010011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0000111010011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0000111010011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000111010011101010) && ({row_reg, col_reg}<19'b0000111010011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000111010011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0000111010011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000111010011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000111010011101111) && ({row_reg, col_reg}<19'b0000111010100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000111010100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0000111010100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0000111010100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0000111010100000100) && ({row_reg, col_reg}<19'b0000111010101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0000111010101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0000111010101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000111010110000000) && ({row_reg, col_reg}<19'b0000111010110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000111010110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0000111010110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0000111010110011010) && ({row_reg, col_reg}<19'b0000111100011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0000111100011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0000111100011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000111100011101010) && ({row_reg, col_reg}<19'b0000111100011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000111100011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0000111100011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000111100011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000111100011101111) && ({row_reg, col_reg}<19'b0000111100100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000111100100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0000111100100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0000111100100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0000111100100000100) && ({row_reg, col_reg}<19'b0000111100101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0000111100101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0000111100101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000111100110000000) && ({row_reg, col_reg}<19'b0000111100110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000111100110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0000111100110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0000111100110011010) && ({row_reg, col_reg}<19'b0000111110011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0000111110011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0000111110011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000111110011101010) && ({row_reg, col_reg}<19'b0000111110011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000111110011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0000111110011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000111110011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000111110011101111) && ({row_reg, col_reg}<19'b0000111110100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000111110100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0000111110100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0000111110100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0000111110100000100) && ({row_reg, col_reg}<19'b0000111110101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0000111110101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0000111110101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000111110110000000) && ({row_reg, col_reg}<19'b0000111110110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000111110110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0000111110110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0000111110110011010) && ({row_reg, col_reg}<19'b0001000000011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0001000000011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0001000000011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0001000000011101010) && ({row_reg, col_reg}<19'b0001000000011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001000000011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0001000000011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001000000011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0001000000011101111) && ({row_reg, col_reg}<19'b0001000000100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001000000100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0001000000100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0001000000100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0001000000100000100) && ({row_reg, col_reg}<19'b0001000000101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0001000000101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0001000000101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0001000000110000000) && ({row_reg, col_reg}<19'b0001000000110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001000000110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0001000000110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0001000000110011010) && ({row_reg, col_reg}<19'b0001000010011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0001000010011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0001000010011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0001000010011101010) && ({row_reg, col_reg}<19'b0001000010011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001000010011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0001000010011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001000010011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0001000010011101111) && ({row_reg, col_reg}<19'b0001000010100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001000010100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0001000010100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0001000010100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0001000010100000100) && ({row_reg, col_reg}<19'b0001000010101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0001000010101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0001000010101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0001000010110000000) && ({row_reg, col_reg}<19'b0001000010110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001000010110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0001000010110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0001000010110011010) && ({row_reg, col_reg}<19'b0001000100011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0001000100011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0001000100011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0001000100011101010) && ({row_reg, col_reg}<19'b0001000100011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001000100011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0001000100011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001000100011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0001000100011101111) && ({row_reg, col_reg}<19'b0001000100100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001000100100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0001000100100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0001000100100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0001000100100000100) && ({row_reg, col_reg}<19'b0001000100101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0001000100101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0001000100101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0001000100110000000) && ({row_reg, col_reg}<19'b0001000100110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001000100110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0001000100110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0001000100110011010) && ({row_reg, col_reg}<19'b0001000110011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0001000110011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0001000110011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0001000110011101010) && ({row_reg, col_reg}<19'b0001000110011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001000110011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0001000110011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001000110011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0001000110011101111) && ({row_reg, col_reg}<19'b0001000110100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001000110100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0001000110100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0001000110100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0001000110100000100) && ({row_reg, col_reg}<19'b0001000110101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0001000110101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0001000110101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0001000110110000000) && ({row_reg, col_reg}<19'b0001000110110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001000110110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0001000110110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0001000110110011010) && ({row_reg, col_reg}<19'b0001001000011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0001001000011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0001001000011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0001001000011101010) && ({row_reg, col_reg}<19'b0001001000011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001001000011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0001001000011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001001000011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0001001000011101111) && ({row_reg, col_reg}<19'b0001001000100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001001000100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0001001000100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0001001000100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0001001000100000100) && ({row_reg, col_reg}<19'b0001001000101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0001001000101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0001001000101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0001001000110000000) && ({row_reg, col_reg}<19'b0001001000110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001001000110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0001001000110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0001001000110011010) && ({row_reg, col_reg}<19'b0001001010011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0001001010011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0001001010011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0001001010011101010) && ({row_reg, col_reg}<19'b0001001010011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001001010011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0001001010011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001001010011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0001001010011101111) && ({row_reg, col_reg}<19'b0001001010100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001001010100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0001001010100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0001001010100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0001001010100000100) && ({row_reg, col_reg}<19'b0001001010101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0001001010101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0001001010101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0001001010110000000) && ({row_reg, col_reg}<19'b0001001010110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001001010110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0001001010110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0001001010110011010) && ({row_reg, col_reg}<19'b0001001100011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0001001100011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0001001100011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0001001100011101010) && ({row_reg, col_reg}<19'b0001001100011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001001100011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0001001100011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001001100011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0001001100011101111) && ({row_reg, col_reg}<19'b0001001100100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001001100100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0001001100100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0001001100100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0001001100100000100) && ({row_reg, col_reg}<19'b0001001100101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0001001100101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0001001100101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0001001100110000000) && ({row_reg, col_reg}<19'b0001001100110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001001100110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0001001100110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0001001100110011010) && ({row_reg, col_reg}<19'b0001001110011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0001001110011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0001001110011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0001001110011101010) && ({row_reg, col_reg}<19'b0001001110011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001001110011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0001001110011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001001110011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0001001110011101111) && ({row_reg, col_reg}<19'b0001001110100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001001110100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0001001110100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0001001110100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0001001110100000100) && ({row_reg, col_reg}<19'b0001001110101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0001001110101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0001001110101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0001001110110000000) && ({row_reg, col_reg}<19'b0001001110110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001001110110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0001001110110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0001001110110011010) && ({row_reg, col_reg}<19'b0001010000011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0001010000011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0001010000011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0001010000011101010) && ({row_reg, col_reg}<19'b0001010000011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001010000011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0001010000011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001010000011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0001010000011101111) && ({row_reg, col_reg}<19'b0001010000100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001010000100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0001010000100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0001010000100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0001010000100000100) && ({row_reg, col_reg}<19'b0001010000101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0001010000101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0001010000101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0001010000110000000) && ({row_reg, col_reg}<19'b0001010000110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001010000110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0001010000110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0001010000110011010) && ({row_reg, col_reg}<19'b0001010010011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0001010010011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0001010010011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0001010010011101010) && ({row_reg, col_reg}<19'b0001010010011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001010010011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0001010010011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001010010011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0001010010011101111) && ({row_reg, col_reg}<19'b0001010010100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001010010100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0001010010100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0001010010100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0001010010100000100) && ({row_reg, col_reg}<19'b0001010010101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0001010010101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0001010010101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0001010010110000000) && ({row_reg, col_reg}<19'b0001010010110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001010010110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0001010010110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0001010010110011010) && ({row_reg, col_reg}<19'b0001010100011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0001010100011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0001010100011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0001010100011101010) && ({row_reg, col_reg}<19'b0001010100011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001010100011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0001010100011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001010100011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0001010100011101111) && ({row_reg, col_reg}<19'b0001010100100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001010100100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0001010100100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0001010100100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0001010100100000100) && ({row_reg, col_reg}<19'b0001010100101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0001010100101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0001010100101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0001010100110000000) && ({row_reg, col_reg}<19'b0001010100110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001010100110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0001010100110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0001010100110011010) && ({row_reg, col_reg}<19'b0001010110011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0001010110011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0001010110011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0001010110011101010) && ({row_reg, col_reg}<19'b0001010110011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001010110011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0001010110011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001010110011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0001010110011101111) && ({row_reg, col_reg}<19'b0001010110100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001010110100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0001010110100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0001010110100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0001010110100000100) && ({row_reg, col_reg}<19'b0001010110101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0001010110101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0001010110101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0001010110110000000) && ({row_reg, col_reg}<19'b0001010110110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001010110110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0001010110110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0001010110110011010) && ({row_reg, col_reg}<19'b0001011000011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0001011000011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0001011000011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0001011000011101010) && ({row_reg, col_reg}<19'b0001011000011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001011000011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0001011000011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001011000011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0001011000011101111) && ({row_reg, col_reg}<19'b0001011000100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001011000100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0001011000100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0001011000100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0001011000100000100) && ({row_reg, col_reg}<19'b0001011000101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0001011000101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0001011000101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0001011000110000000) && ({row_reg, col_reg}<19'b0001011000110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001011000110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0001011000110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0001011000110011010) && ({row_reg, col_reg}<19'b0001011010011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0001011010011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0001011010011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0001011010011101010) && ({row_reg, col_reg}<19'b0001011010011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001011010011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0001011010011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001011010011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0001011010011101111) && ({row_reg, col_reg}<19'b0001011010100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001011010100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0001011010100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0001011010100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0001011010100000100) && ({row_reg, col_reg}<19'b0001011010101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0001011010101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0001011010101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0001011010110000000) && ({row_reg, col_reg}<19'b0001011010110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001011010110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0001011010110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0001011010110011010) && ({row_reg, col_reg}<19'b0001011100011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0001011100011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0001011100011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0001011100011101010) && ({row_reg, col_reg}<19'b0001011100011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001011100011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0001011100011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001011100011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0001011100011101111) && ({row_reg, col_reg}<19'b0001011100100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001011100100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0001011100100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0001011100100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0001011100100000100) && ({row_reg, col_reg}<19'b0001011100101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0001011100101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0001011100101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0001011100110000000) && ({row_reg, col_reg}<19'b0001011100110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001011100110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0001011100110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0001011100110011010) && ({row_reg, col_reg}<19'b0001011110011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0001011110011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0001011110011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0001011110011101010) && ({row_reg, col_reg}<19'b0001011110011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001011110011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0001011110011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001011110011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0001011110011101111) && ({row_reg, col_reg}<19'b0001011110100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001011110100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0001011110100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0001011110100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0001011110100000100) && ({row_reg, col_reg}<19'b0001011110101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0001011110101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0001011110101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0001011110110000000) && ({row_reg, col_reg}<19'b0001011110110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001011110110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0001011110110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0001011110110011010) && ({row_reg, col_reg}<19'b0001100000011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0001100000011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0001100000011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0001100000011101010) && ({row_reg, col_reg}<19'b0001100000011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001100000011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0001100000011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001100000011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0001100000011101111) && ({row_reg, col_reg}<19'b0001100000100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001100000100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0001100000100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0001100000100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0001100000100000100) && ({row_reg, col_reg}<19'b0001100000101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0001100000101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0001100000101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0001100000110000000) && ({row_reg, col_reg}<19'b0001100000110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001100000110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0001100000110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0001100000110011010) && ({row_reg, col_reg}<19'b0001100010011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0001100010011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0001100010011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0001100010011101010) && ({row_reg, col_reg}<19'b0001100010011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001100010011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0001100010011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001100010011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0001100010011101111) && ({row_reg, col_reg}<19'b0001100010100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001100010100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0001100010100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0001100010100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0001100010100000100) && ({row_reg, col_reg}<19'b0001100010101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0001100010101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0001100010101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0001100010110000000) && ({row_reg, col_reg}<19'b0001100010110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001100010110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0001100010110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0001100010110011010) && ({row_reg, col_reg}<19'b0001100100011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0001100100011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0001100100011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0001100100011101010) && ({row_reg, col_reg}<19'b0001100100011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001100100011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0001100100011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001100100011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0001100100011101111) && ({row_reg, col_reg}<19'b0001100100100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001100100100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0001100100100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0001100100100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0001100100100000100) && ({row_reg, col_reg}<19'b0001100100101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0001100100101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0001100100101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0001100100110000000) && ({row_reg, col_reg}<19'b0001100100110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001100100110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0001100100110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0001100100110011010) && ({row_reg, col_reg}<19'b0001100110011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0001100110011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0001100110011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0001100110011101010) && ({row_reg, col_reg}<19'b0001100110011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001100110011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0001100110011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001100110011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0001100110011101111) && ({row_reg, col_reg}<19'b0001100110100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001100110100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0001100110100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0001100110100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0001100110100000100) && ({row_reg, col_reg}<19'b0001100110101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0001100110101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0001100110101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0001100110110000000) && ({row_reg, col_reg}<19'b0001100110110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001100110110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0001100110110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0001100110110011010) && ({row_reg, col_reg}<19'b0001101000011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0001101000011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0001101000011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0001101000011101010) && ({row_reg, col_reg}<19'b0001101000011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001101000011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0001101000011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001101000011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0001101000011101111) && ({row_reg, col_reg}<19'b0001101000100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001101000100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0001101000100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0001101000100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0001101000100000100) && ({row_reg, col_reg}<19'b0001101000101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0001101000101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0001101000101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0001101000110000000) && ({row_reg, col_reg}<19'b0001101000110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001101000110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0001101000110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0001101000110011010) && ({row_reg, col_reg}<19'b0001101010011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0001101010011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0001101010011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0001101010011101010) && ({row_reg, col_reg}<19'b0001101010011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001101010011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0001101010011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001101010011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0001101010011101111) && ({row_reg, col_reg}<19'b0001101010100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001101010100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0001101010100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0001101010100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0001101010100000100) && ({row_reg, col_reg}<19'b0001101010101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0001101010101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0001101010101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0001101010110000000) && ({row_reg, col_reg}<19'b0001101010110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001101010110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0001101010110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0001101010110011010) && ({row_reg, col_reg}<19'b0001101100011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0001101100011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0001101100011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0001101100011101010) && ({row_reg, col_reg}<19'b0001101100011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001101100011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0001101100011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001101100011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0001101100011101111) && ({row_reg, col_reg}<19'b0001101100100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001101100100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0001101100100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0001101100100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0001101100100000100) && ({row_reg, col_reg}<19'b0001101100101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0001101100101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0001101100101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0001101100110000000) && ({row_reg, col_reg}<19'b0001101100110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001101100110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0001101100110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0001101100110011010) && ({row_reg, col_reg}<19'b0001101110011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0001101110011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0001101110011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0001101110011101010) && ({row_reg, col_reg}<19'b0001101110011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001101110011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0001101110011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001101110011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0001101110011101111) && ({row_reg, col_reg}<19'b0001101110100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001101110100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0001101110100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0001101110100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0001101110100000100) && ({row_reg, col_reg}<19'b0001101110101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0001101110101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0001101110101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0001101110110000000) && ({row_reg, col_reg}<19'b0001101110110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001101110110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0001101110110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0001101110110011010) && ({row_reg, col_reg}<19'b0001110000011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0001110000011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0001110000011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0001110000011101010) && ({row_reg, col_reg}<19'b0001110000011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001110000011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0001110000011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001110000011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0001110000011101111) && ({row_reg, col_reg}<19'b0001110000100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001110000100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0001110000100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0001110000100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0001110000100000100) && ({row_reg, col_reg}<19'b0001110000101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0001110000101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0001110000101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0001110000110000000) && ({row_reg, col_reg}<19'b0001110000110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001110000110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0001110000110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0001110000110011010) && ({row_reg, col_reg}<19'b0001110010011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0001110010011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0001110010011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0001110010011101010) && ({row_reg, col_reg}<19'b0001110010011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001110010011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0001110010011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001110010011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0001110010011101111) && ({row_reg, col_reg}<19'b0001110010100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001110010100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0001110010100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0001110010100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0001110010100000100) && ({row_reg, col_reg}<19'b0001110010101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0001110010101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0001110010101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0001110010110000000) && ({row_reg, col_reg}<19'b0001110010110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001110010110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0001110010110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0001110010110011010) && ({row_reg, col_reg}<19'b0001110100011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0001110100011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0001110100011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0001110100011101010) && ({row_reg, col_reg}<19'b0001110100011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001110100011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0001110100011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001110100011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0001110100011101111) && ({row_reg, col_reg}<19'b0001110100100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001110100100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0001110100100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0001110100100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0001110100100000100) && ({row_reg, col_reg}<19'b0001110100101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0001110100101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0001110100101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0001110100110000000) && ({row_reg, col_reg}<19'b0001110100110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001110100110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0001110100110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0001110100110011010) && ({row_reg, col_reg}<19'b0001110110011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0001110110011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0001110110011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0001110110011101010) && ({row_reg, col_reg}<19'b0001110110011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001110110011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0001110110011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001110110011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0001110110011101111) && ({row_reg, col_reg}<19'b0001110110100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001110110100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0001110110100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0001110110100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0001110110100000100) && ({row_reg, col_reg}<19'b0001110110101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0001110110101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0001110110101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0001110110110000000) && ({row_reg, col_reg}<19'b0001110110110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001110110110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0001110110110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0001110110110011010) && ({row_reg, col_reg}<19'b0001111000011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0001111000011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0001111000011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0001111000011101010) && ({row_reg, col_reg}<19'b0001111000011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001111000011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0001111000011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001111000011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0001111000011101111) && ({row_reg, col_reg}<19'b0001111000100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001111000100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0001111000100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0001111000100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0001111000100000100) && ({row_reg, col_reg}<19'b0001111000101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0001111000101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0001111000101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0001111000110000000) && ({row_reg, col_reg}<19'b0001111000110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001111000110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0001111000110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0001111000110011010) && ({row_reg, col_reg}<19'b0001111010011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0001111010011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0001111010011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0001111010011101010) && ({row_reg, col_reg}<19'b0001111010011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001111010011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0001111010011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001111010011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0001111010011101111) && ({row_reg, col_reg}<19'b0001111010100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001111010100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0001111010100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0001111010100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0001111010100000100) && ({row_reg, col_reg}<19'b0001111010101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0001111010101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0001111010101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0001111010110000000) && ({row_reg, col_reg}<19'b0001111010110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001111010110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0001111010110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0001111010110011010) && ({row_reg, col_reg}<19'b0001111100011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0001111100011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0001111100011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0001111100011101010) && ({row_reg, col_reg}<19'b0001111100011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001111100011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0001111100011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001111100011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0001111100011101111) && ({row_reg, col_reg}<19'b0001111100100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001111100100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0001111100100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0001111100100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0001111100100000100) && ({row_reg, col_reg}<19'b0001111100101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0001111100101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0001111100101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0001111100110000000) && ({row_reg, col_reg}<19'b0001111100110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001111100110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0001111100110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0001111100110011010) && ({row_reg, col_reg}<19'b0001111110011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0001111110011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0001111110011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0001111110011101010) && ({row_reg, col_reg}<19'b0001111110011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001111110011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0001111110011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001111110011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0001111110011101111) && ({row_reg, col_reg}<19'b0001111110100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001111110100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0001111110100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0001111110100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0001111110100000100) && ({row_reg, col_reg}<19'b0001111110101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0001111110101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0001111110101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0001111110110000000) && ({row_reg, col_reg}<19'b0001111110110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001111110110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0001111110110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0001111110110011010) && ({row_reg, col_reg}<19'b0010000000011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010000000011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0010000000011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010000000011101010) && ({row_reg, col_reg}<19'b0010000000011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010000000011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0010000000011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010000000011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010000000011101111) && ({row_reg, col_reg}<19'b0010000000100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010000000100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0010000000100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0010000000100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0010000000100000100) && ({row_reg, col_reg}<19'b0010000000101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010000000101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0010000000101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010000000110000000) && ({row_reg, col_reg}<19'b0010000000110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010000000110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0010000000110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0010000000110011010) && ({row_reg, col_reg}<19'b0010000010011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010000010011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0010000010011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010000010011101010) && ({row_reg, col_reg}<19'b0010000010011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010000010011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0010000010011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010000010011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010000010011101111) && ({row_reg, col_reg}<19'b0010000010100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010000010100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0010000010100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0010000010100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0010000010100000100) && ({row_reg, col_reg}<19'b0010000010101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010000010101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0010000010101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010000010110000000) && ({row_reg, col_reg}<19'b0010000010110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010000010110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0010000010110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0010000010110011010) && ({row_reg, col_reg}<19'b0010000100011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010000100011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0010000100011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010000100011101010) && ({row_reg, col_reg}<19'b0010000100011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010000100011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0010000100011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010000100011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010000100011101111) && ({row_reg, col_reg}<19'b0010000100100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010000100100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0010000100100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0010000100100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0010000100100000100) && ({row_reg, col_reg}<19'b0010000100101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010000100101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0010000100101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010000100110000000) && ({row_reg, col_reg}<19'b0010000100110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010000100110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0010000100110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0010000100110011010) && ({row_reg, col_reg}<19'b0010000110011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010000110011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0010000110011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010000110011101010) && ({row_reg, col_reg}<19'b0010000110011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010000110011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0010000110011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010000110011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010000110011101111) && ({row_reg, col_reg}<19'b0010000110100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010000110100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0010000110100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0010000110100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0010000110100000100) && ({row_reg, col_reg}<19'b0010000110101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010000110101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0010000110101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010000110110000000) && ({row_reg, col_reg}<19'b0010000110110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010000110110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0010000110110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0010000110110011010) && ({row_reg, col_reg}<19'b0010001000011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010001000011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0010001000011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010001000011101010) && ({row_reg, col_reg}<19'b0010001000011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010001000011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0010001000011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010001000011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010001000011101111) && ({row_reg, col_reg}<19'b0010001000100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010001000100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0010001000100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0010001000100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0010001000100000100) && ({row_reg, col_reg}<19'b0010001000101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010001000101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0010001000101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010001000110000000) && ({row_reg, col_reg}<19'b0010001000110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010001000110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0010001000110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0010001000110011010) && ({row_reg, col_reg}<19'b0010001010011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010001010011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0010001010011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010001010011101010) && ({row_reg, col_reg}<19'b0010001010011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010001010011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0010001010011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010001010011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010001010011101111) && ({row_reg, col_reg}<19'b0010001010100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010001010100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0010001010100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0010001010100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0010001010100000100) && ({row_reg, col_reg}<19'b0010001010101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010001010101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0010001010101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010001010110000000) && ({row_reg, col_reg}<19'b0010001010110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010001010110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0010001010110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0010001010110011010) && ({row_reg, col_reg}<19'b0010001100011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010001100011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0010001100011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010001100011101010) && ({row_reg, col_reg}<19'b0010001100011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010001100011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0010001100011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010001100011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010001100011101111) && ({row_reg, col_reg}<19'b0010001100100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010001100100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0010001100100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0010001100100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0010001100100000100) && ({row_reg, col_reg}<19'b0010001100101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010001100101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0010001100101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010001100110000000) && ({row_reg, col_reg}<19'b0010001100110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010001100110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0010001100110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0010001100110011010) && ({row_reg, col_reg}<19'b0010001110011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010001110011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0010001110011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010001110011101010) && ({row_reg, col_reg}<19'b0010001110011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010001110011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0010001110011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010001110011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010001110011101111) && ({row_reg, col_reg}<19'b0010001110100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010001110100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0010001110100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0010001110100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0010001110100000100) && ({row_reg, col_reg}<19'b0010001110101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010001110101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0010001110101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010001110110000000) && ({row_reg, col_reg}<19'b0010001110110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010001110110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0010001110110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0010001110110011010) && ({row_reg, col_reg}<19'b0010010000011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010010000011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0010010000011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010010000011101010) && ({row_reg, col_reg}<19'b0010010000011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010010000011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0010010000011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010010000011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010010000011101111) && ({row_reg, col_reg}<19'b0010010000100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010010000100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0010010000100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0010010000100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0010010000100000100) && ({row_reg, col_reg}<19'b0010010000101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010010000101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0010010000101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010010000110000000) && ({row_reg, col_reg}<19'b0010010000110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010010000110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0010010000110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0010010000110011010) && ({row_reg, col_reg}<19'b0010010010011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010010010011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0010010010011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010010010011101010) && ({row_reg, col_reg}<19'b0010010010011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010010010011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0010010010011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010010010011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010010010011101111) && ({row_reg, col_reg}<19'b0010010010100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010010010100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0010010010100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0010010010100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0010010010100000100) && ({row_reg, col_reg}<19'b0010010010101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010010010101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0010010010101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010010010110000000) && ({row_reg, col_reg}<19'b0010010010110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010010010110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0010010010110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0010010010110011010) && ({row_reg, col_reg}<19'b0010010100011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010010100011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0010010100011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010010100011101010) && ({row_reg, col_reg}<19'b0010010100011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010010100011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0010010100011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010010100011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010010100011101111) && ({row_reg, col_reg}<19'b0010010100100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010010100100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0010010100100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0010010100100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0010010100100000100) && ({row_reg, col_reg}<19'b0010010100101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010010100101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0010010100101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010010100110000000) && ({row_reg, col_reg}<19'b0010010100110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010010100110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0010010100110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0010010100110011010) && ({row_reg, col_reg}<19'b0010010110011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010010110011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0010010110011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010010110011101010) && ({row_reg, col_reg}<19'b0010010110011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010010110011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0010010110011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010010110011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010010110011101111) && ({row_reg, col_reg}<19'b0010010110100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010010110100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0010010110100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0010010110100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0010010110100000100) && ({row_reg, col_reg}<19'b0010010110101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010010110101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0010010110101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010010110110000000) && ({row_reg, col_reg}<19'b0010010110110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010010110110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0010010110110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0010010110110011010) && ({row_reg, col_reg}<19'b0010011000011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010011000011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0010011000011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010011000011101010) && ({row_reg, col_reg}<19'b0010011000011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010011000011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0010011000011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010011000011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010011000011101111) && ({row_reg, col_reg}<19'b0010011000100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010011000100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0010011000100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0010011000100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0010011000100000100) && ({row_reg, col_reg}<19'b0010011000101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010011000101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0010011000101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010011000110000000) && ({row_reg, col_reg}<19'b0010011000110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010011000110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0010011000110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0010011000110011010) && ({row_reg, col_reg}<19'b0010011010011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010011010011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0010011010011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010011010011101010) && ({row_reg, col_reg}<19'b0010011010011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010011010011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0010011010011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010011010011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010011010011101111) && ({row_reg, col_reg}<19'b0010011010100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010011010100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0010011010100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0010011010100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0010011010100000100) && ({row_reg, col_reg}<19'b0010011010101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010011010101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0010011010101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010011010110000000) && ({row_reg, col_reg}<19'b0010011010110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010011010110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0010011010110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0010011010110011010) && ({row_reg, col_reg}<19'b0010011100011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010011100011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0010011100011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010011100011101010) && ({row_reg, col_reg}<19'b0010011100011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010011100011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0010011100011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010011100011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010011100011101111) && ({row_reg, col_reg}<19'b0010011100100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010011100100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0010011100100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0010011100100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0010011100100000100) && ({row_reg, col_reg}<19'b0010011100101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010011100101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0010011100101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010011100110000000) && ({row_reg, col_reg}<19'b0010011100110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010011100110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0010011100110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0010011100110011010) && ({row_reg, col_reg}<19'b0010011110011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010011110011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0010011110011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010011110011101010) && ({row_reg, col_reg}<19'b0010011110011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010011110011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0010011110011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010011110011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010011110011101111) && ({row_reg, col_reg}<19'b0010011110100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010011110100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0010011110100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0010011110100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0010011110100000100) && ({row_reg, col_reg}<19'b0010011110101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010011110101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0010011110101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010011110110000000) && ({row_reg, col_reg}<19'b0010011110110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010011110110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0010011110110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0010011110110011010) && ({row_reg, col_reg}<19'b0010100000011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010100000011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0010100000011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010100000011101010) && ({row_reg, col_reg}<19'b0010100000011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010100000011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0010100000011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010100000011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010100000011101111) && ({row_reg, col_reg}<19'b0010100000100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010100000100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0010100000100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0010100000100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0010100000100000100) && ({row_reg, col_reg}<19'b0010100000101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010100000101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0010100000101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010100000110000000) && ({row_reg, col_reg}<19'b0010100000110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010100000110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0010100000110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0010100000110011010) && ({row_reg, col_reg}<19'b0010100010011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010100010011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0010100010011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010100010011101010) && ({row_reg, col_reg}<19'b0010100010011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010100010011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0010100010011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010100010011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010100010011101111) && ({row_reg, col_reg}<19'b0010100010100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010100010100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0010100010100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0010100010100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0010100010100000100) && ({row_reg, col_reg}<19'b0010100010101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010100010101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0010100010101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010100010110000000) && ({row_reg, col_reg}<19'b0010100010110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010100010110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0010100010110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0010100010110011010) && ({row_reg, col_reg}<19'b0010100100011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010100100011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0010100100011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010100100011101010) && ({row_reg, col_reg}<19'b0010100100011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010100100011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0010100100011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010100100011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010100100011101111) && ({row_reg, col_reg}<19'b0010100100100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010100100100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0010100100100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0010100100100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0010100100100000100) && ({row_reg, col_reg}<19'b0010100100101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010100100101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0010100100101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010100100110000000) && ({row_reg, col_reg}<19'b0010100100110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010100100110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0010100100110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0010100100110011010) && ({row_reg, col_reg}<19'b0010100110011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010100110011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0010100110011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010100110011101010) && ({row_reg, col_reg}<19'b0010100110011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010100110011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0010100110011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010100110011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010100110011101111) && ({row_reg, col_reg}<19'b0010100110100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010100110100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0010100110100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0010100110100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0010100110100000100) && ({row_reg, col_reg}<19'b0010100110101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010100110101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0010100110101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010100110110000000) && ({row_reg, col_reg}<19'b0010100110110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010100110110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0010100110110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0010100110110011010) && ({row_reg, col_reg}<19'b0010101000011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010101000011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0010101000011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010101000011101010) && ({row_reg, col_reg}<19'b0010101000011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010101000011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0010101000011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010101000011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010101000011101111) && ({row_reg, col_reg}<19'b0010101000100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010101000100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0010101000100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0010101000100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0010101000100000100) && ({row_reg, col_reg}<19'b0010101000101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010101000101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0010101000101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010101000110000000) && ({row_reg, col_reg}<19'b0010101000110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010101000110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0010101000110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0010101000110011010) && ({row_reg, col_reg}<19'b0010101010011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010101010011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0010101010011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010101010011101010) && ({row_reg, col_reg}<19'b0010101010011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010101010011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0010101010011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010101010011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010101010011101111) && ({row_reg, col_reg}<19'b0010101010100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010101010100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0010101010100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0010101010100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0010101010100000100) && ({row_reg, col_reg}<19'b0010101010101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010101010101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0010101010101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010101010110000000) && ({row_reg, col_reg}<19'b0010101010110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010101010110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0010101010110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0010101010110011010) && ({row_reg, col_reg}<19'b0010101100011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010101100011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0010101100011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010101100011101010) && ({row_reg, col_reg}<19'b0010101100011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010101100011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0010101100011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010101100011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010101100011101111) && ({row_reg, col_reg}<19'b0010101100100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010101100100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0010101100100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0010101100100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0010101100100000100) && ({row_reg, col_reg}<19'b0010101100101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010101100101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0010101100101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010101100110000000) && ({row_reg, col_reg}<19'b0010101100110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010101100110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0010101100110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0010101100110011010) && ({row_reg, col_reg}<19'b0010101110011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010101110011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0010101110011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010101110011101010) && ({row_reg, col_reg}<19'b0010101110011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010101110011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0010101110011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010101110011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010101110011101111) && ({row_reg, col_reg}<19'b0010101110100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010101110100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0010101110100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0010101110100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0010101110100000100) && ({row_reg, col_reg}<19'b0010101110101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010101110101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0010101110101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010101110110000000) && ({row_reg, col_reg}<19'b0010101110110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010101110110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0010101110110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0010101110110011010) && ({row_reg, col_reg}<19'b0010110000011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010110000011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0010110000011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010110000011101010) && ({row_reg, col_reg}<19'b0010110000011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010110000011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0010110000011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010110000011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010110000011101111) && ({row_reg, col_reg}<19'b0010110000100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010110000100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0010110000100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0010110000100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0010110000100000100) && ({row_reg, col_reg}<19'b0010110000101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010110000101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0010110000101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010110000110000000) && ({row_reg, col_reg}<19'b0010110000110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010110000110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0010110000110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0010110000110011010) && ({row_reg, col_reg}<19'b0010110010011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010110010011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0010110010011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010110010011101010) && ({row_reg, col_reg}<19'b0010110010011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010110010011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0010110010011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010110010011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010110010011101111) && ({row_reg, col_reg}<19'b0010110010100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010110010100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0010110010100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0010110010100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0010110010100000100) && ({row_reg, col_reg}<19'b0010110010101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010110010101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0010110010101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010110010110000000) && ({row_reg, col_reg}<19'b0010110010110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010110010110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0010110010110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0010110010110011010) && ({row_reg, col_reg}<19'b0010110100011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010110100011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0010110100011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010110100011101010) && ({row_reg, col_reg}<19'b0010110100011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010110100011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0010110100011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010110100011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010110100011101111) && ({row_reg, col_reg}<19'b0010110100100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010110100100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0010110100100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0010110100100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0010110100100000100) && ({row_reg, col_reg}<19'b0010110100101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010110100101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0010110100101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010110100110000000) && ({row_reg, col_reg}<19'b0010110100110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010110100110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0010110100110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0010110100110011010) && ({row_reg, col_reg}<19'b0010110110011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010110110011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0010110110011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010110110011101010) && ({row_reg, col_reg}<19'b0010110110011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010110110011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0010110110011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010110110011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010110110011101111) && ({row_reg, col_reg}<19'b0010110110100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010110110100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0010110110100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0010110110100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0010110110100000100) && ({row_reg, col_reg}<19'b0010110110101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010110110101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0010110110101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010110110110000000) && ({row_reg, col_reg}<19'b0010110110110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010110110110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0010110110110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0010110110110011010) && ({row_reg, col_reg}<19'b0010111000011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010111000011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0010111000011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010111000011101010) && ({row_reg, col_reg}<19'b0010111000011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010111000011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0010111000011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010111000011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010111000011101111) && ({row_reg, col_reg}<19'b0010111000100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010111000100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0010111000100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0010111000100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0010111000100000100) && ({row_reg, col_reg}<19'b0010111000101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010111000101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0010111000101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010111000110000000) && ({row_reg, col_reg}<19'b0010111000110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010111000110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0010111000110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0010111000110011010) && ({row_reg, col_reg}<19'b0010111010011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010111010011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0010111010011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010111010011101010) && ({row_reg, col_reg}<19'b0010111010011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010111010011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0010111010011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010111010011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010111010011101111) && ({row_reg, col_reg}<19'b0010111010100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010111010100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0010111010100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0010111010100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0010111010100000100) && ({row_reg, col_reg}<19'b0010111010101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010111010101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0010111010101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010111010110000000) && ({row_reg, col_reg}<19'b0010111010110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010111010110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0010111010110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0010111010110011010) && ({row_reg, col_reg}<19'b0010111100011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010111100011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0010111100011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010111100011101010) && ({row_reg, col_reg}<19'b0010111100011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010111100011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0010111100011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010111100011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010111100011101111) && ({row_reg, col_reg}<19'b0010111100100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010111100100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0010111100100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0010111100100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0010111100100000100) && ({row_reg, col_reg}<19'b0010111100101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010111100101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0010111100101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010111100110000000) && ({row_reg, col_reg}<19'b0010111100110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010111100110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0010111100110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0010111100110011010) && ({row_reg, col_reg}<19'b0010111110011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010111110011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0010111110011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010111110011101010) && ({row_reg, col_reg}<19'b0010111110011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010111110011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0010111110011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010111110011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010111110011101111) && ({row_reg, col_reg}<19'b0010111110100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010111110100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0010111110100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0010111110100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0010111110100000100) && ({row_reg, col_reg}<19'b0010111110101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010111110101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0010111110101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010111110110000000) && ({row_reg, col_reg}<19'b0010111110110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010111110110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0010111110110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0010111110110011010) && ({row_reg, col_reg}<19'b0011000000011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011000000011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0011000000011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011000000011101010) && ({row_reg, col_reg}<19'b0011000000011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011000000011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011000000011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011000000011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011000000011101111) && ({row_reg, col_reg}<19'b0011000000100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011000000100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011000000100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0011000000100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0011000000100000100) && ({row_reg, col_reg}<19'b0011000000101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011000000101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0011000000101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011000000110000000) && ({row_reg, col_reg}<19'b0011000000110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011000000110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0011000000110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0011000000110011010) && ({row_reg, col_reg}<19'b0011000010011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011000010011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0011000010011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011000010011101010) && ({row_reg, col_reg}<19'b0011000010011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011000010011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011000010011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011000010011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011000010011101111) && ({row_reg, col_reg}<19'b0011000010100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011000010100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011000010100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0011000010100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0011000010100000100) && ({row_reg, col_reg}<19'b0011000010101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011000010101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0011000010101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011000010110000000) && ({row_reg, col_reg}<19'b0011000010110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011000010110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0011000010110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0011000010110011010) && ({row_reg, col_reg}<19'b0011000100011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011000100011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0011000100011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011000100011101010) && ({row_reg, col_reg}<19'b0011000100011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011000100011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011000100011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011000100011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011000100011101111) && ({row_reg, col_reg}<19'b0011000100100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011000100100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011000100100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0011000100100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0011000100100000100) && ({row_reg, col_reg}<19'b0011000100101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011000100101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0011000100101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011000100110000000) && ({row_reg, col_reg}<19'b0011000100110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011000100110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0011000100110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0011000100110011010) && ({row_reg, col_reg}<19'b0011000110011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011000110011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0011000110011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011000110011101010) && ({row_reg, col_reg}<19'b0011000110011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011000110011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011000110011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011000110011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011000110011101111) && ({row_reg, col_reg}<19'b0011000110100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011000110100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011000110100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0011000110100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0011000110100000100) && ({row_reg, col_reg}<19'b0011000110101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011000110101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0011000110101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011000110110000000) && ({row_reg, col_reg}<19'b0011000110110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011000110110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0011000110110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0011000110110011010) && ({row_reg, col_reg}<19'b0011001000011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011001000011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0011001000011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011001000011101010) && ({row_reg, col_reg}<19'b0011001000011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011001000011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011001000011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011001000011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011001000011101111) && ({row_reg, col_reg}<19'b0011001000100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011001000100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011001000100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0011001000100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0011001000100000100) && ({row_reg, col_reg}<19'b0011001000101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011001000101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0011001000101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011001000110000000) && ({row_reg, col_reg}<19'b0011001000110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011001000110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0011001000110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0011001000110011010) && ({row_reg, col_reg}<19'b0011001010011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011001010011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0011001010011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011001010011101010) && ({row_reg, col_reg}<19'b0011001010011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011001010011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011001010011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011001010011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011001010011101111) && ({row_reg, col_reg}<19'b0011001010100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011001010100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011001010100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0011001010100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0011001010100000100) && ({row_reg, col_reg}<19'b0011001010101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011001010101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0011001010101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011001010110000000) && ({row_reg, col_reg}<19'b0011001010110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011001010110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0011001010110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0011001010110011010) && ({row_reg, col_reg}<19'b0011001100011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011001100011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0011001100011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011001100011101010) && ({row_reg, col_reg}<19'b0011001100011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011001100011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011001100011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011001100011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011001100011101111) && ({row_reg, col_reg}<19'b0011001100100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011001100100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011001100100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0011001100100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0011001100100000100) && ({row_reg, col_reg}<19'b0011001100101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011001100101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0011001100101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011001100110000000) && ({row_reg, col_reg}<19'b0011001100110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011001100110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0011001100110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0011001100110011010) && ({row_reg, col_reg}<19'b0011001110011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011001110011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0011001110011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011001110011101010) && ({row_reg, col_reg}<19'b0011001110011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011001110011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011001110011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011001110011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011001110011101111) && ({row_reg, col_reg}<19'b0011001110100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011001110100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011001110100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0011001110100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0011001110100000100) && ({row_reg, col_reg}<19'b0011001110101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011001110101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0011001110101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011001110110000000) && ({row_reg, col_reg}<19'b0011001110110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011001110110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0011001110110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0011001110110011010) && ({row_reg, col_reg}<19'b0011010000011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011010000011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0011010000011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011010000011101010) && ({row_reg, col_reg}<19'b0011010000011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011010000011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011010000011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011010000011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011010000011101111) && ({row_reg, col_reg}<19'b0011010000100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011010000100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011010000100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0011010000100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0011010000100000100) && ({row_reg, col_reg}<19'b0011010000101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011010000101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0011010000101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011010000110000000) && ({row_reg, col_reg}<19'b0011010000110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011010000110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0011010000110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0011010000110011010) && ({row_reg, col_reg}<19'b0011010010011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011010010011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0011010010011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011010010011101010) && ({row_reg, col_reg}<19'b0011010010011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011010010011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011010010011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011010010011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011010010011101111) && ({row_reg, col_reg}<19'b0011010010100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011010010100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011010010100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0011010010100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0011010010100000100) && ({row_reg, col_reg}<19'b0011010010101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011010010101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0011010010101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011010010110000000) && ({row_reg, col_reg}<19'b0011010010110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011010010110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0011010010110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0011010010110011010) && ({row_reg, col_reg}<19'b0011010100011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011010100011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0011010100011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011010100011101010) && ({row_reg, col_reg}<19'b0011010100011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011010100011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011010100011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011010100011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011010100011101111) && ({row_reg, col_reg}<19'b0011010100100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011010100100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011010100100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0011010100100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0011010100100000100) && ({row_reg, col_reg}<19'b0011010100101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011010100101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0011010100101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011010100110000000) && ({row_reg, col_reg}<19'b0011010100110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011010100110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0011010100110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0011010100110011010) && ({row_reg, col_reg}<19'b0011010110011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011010110011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0011010110011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011010110011101010) && ({row_reg, col_reg}<19'b0011010110011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011010110011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011010110011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011010110011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011010110011101111) && ({row_reg, col_reg}<19'b0011010110100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011010110100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011010110100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0011010110100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0011010110100000100) && ({row_reg, col_reg}<19'b0011010110101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011010110101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0011010110101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011010110110000000) && ({row_reg, col_reg}<19'b0011010110110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011010110110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0011010110110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0011010110110011010) && ({row_reg, col_reg}<19'b0011011000011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011011000011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0011011000011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011011000011101010) && ({row_reg, col_reg}<19'b0011011000011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011011000011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011011000011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011011000011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011011000011101111) && ({row_reg, col_reg}<19'b0011011000100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011011000100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011011000100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0011011000100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0011011000100000100) && ({row_reg, col_reg}<19'b0011011000101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011011000101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0011011000101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011011000110000000) && ({row_reg, col_reg}<19'b0011011000110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011011000110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0011011000110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0011011000110011010) && ({row_reg, col_reg}<19'b0011011010011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011011010011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0011011010011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011011010011101010) && ({row_reg, col_reg}<19'b0011011010011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011011010011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011011010011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011011010011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011011010011101111) && ({row_reg, col_reg}<19'b0011011010100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011011010100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011011010100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0011011010100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0011011010100000100) && ({row_reg, col_reg}<19'b0011011010101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011011010101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0011011010101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011011010110000000) && ({row_reg, col_reg}<19'b0011011010110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011011010110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0011011010110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0011011010110011010) && ({row_reg, col_reg}<19'b0011011100011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011011100011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0011011100011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011011100011101010) && ({row_reg, col_reg}<19'b0011011100011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011011100011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011011100011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011011100011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011011100011101111) && ({row_reg, col_reg}<19'b0011011100100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011011100100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011011100100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0011011100100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0011011100100000100) && ({row_reg, col_reg}<19'b0011011100101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011011100101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0011011100101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011011100110000000) && ({row_reg, col_reg}<19'b0011011100110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011011100110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0011011100110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0011011100110011010) && ({row_reg, col_reg}<19'b0011011110011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011011110011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0011011110011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011011110011101010) && ({row_reg, col_reg}<19'b0011011110011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011011110011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011011110011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011011110011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011011110011101111) && ({row_reg, col_reg}<19'b0011011110100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011011110100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011011110100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0011011110100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0011011110100000100) && ({row_reg, col_reg}<19'b0011011110101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011011110101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0011011110101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011011110110000000) && ({row_reg, col_reg}<19'b0011011110110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011011110110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0011011110110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0011011110110011010) && ({row_reg, col_reg}<19'b0011100000011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011100000011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0011100000011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011100000011101010) && ({row_reg, col_reg}<19'b0011100000011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011100000011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011100000011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011100000011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011100000011101111) && ({row_reg, col_reg}<19'b0011100000100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011100000100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011100000100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0011100000100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0011100000100000100) && ({row_reg, col_reg}<19'b0011100000101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011100000101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0011100000101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011100000110000000) && ({row_reg, col_reg}<19'b0011100000110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011100000110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0011100000110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0011100000110011010) && ({row_reg, col_reg}<19'b0011100010011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011100010011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0011100010011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011100010011101010) && ({row_reg, col_reg}<19'b0011100010011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011100010011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011100010011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011100010011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011100010011101111) && ({row_reg, col_reg}<19'b0011100010100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011100010100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011100010100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0011100010100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0011100010100000100) && ({row_reg, col_reg}<19'b0011100010101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011100010101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0011100010101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011100010110000000) && ({row_reg, col_reg}<19'b0011100010110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011100010110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0011100010110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0011100010110011010) && ({row_reg, col_reg}<19'b0011100100011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011100100011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0011100100011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011100100011101010) && ({row_reg, col_reg}<19'b0011100100011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011100100011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011100100011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011100100011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011100100011101111) && ({row_reg, col_reg}<19'b0011100100100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011100100100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011100100100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0011100100100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0011100100100000100) && ({row_reg, col_reg}<19'b0011100100101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011100100101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0011100100101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011100100110000000) && ({row_reg, col_reg}<19'b0011100100110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011100100110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0011100100110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0011100100110011010) && ({row_reg, col_reg}<19'b0011100110011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011100110011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0011100110011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011100110011101010) && ({row_reg, col_reg}<19'b0011100110011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011100110011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011100110011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011100110011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011100110011101111) && ({row_reg, col_reg}<19'b0011100110100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011100110100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011100110100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0011100110100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0011100110100000100) && ({row_reg, col_reg}<19'b0011100110101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011100110101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0011100110101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011100110110000000) && ({row_reg, col_reg}<19'b0011100110110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011100110110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0011100110110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0011100110110011010) && ({row_reg, col_reg}<19'b0011101000011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011101000011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0011101000011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011101000011101010) && ({row_reg, col_reg}<19'b0011101000011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011101000011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011101000011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011101000011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011101000011101111) && ({row_reg, col_reg}<19'b0011101000100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011101000100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011101000100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0011101000100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0011101000100000100) && ({row_reg, col_reg}<19'b0011101000101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011101000101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0011101000101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011101000110000000) && ({row_reg, col_reg}<19'b0011101000110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011101000110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0011101000110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0011101000110011010) && ({row_reg, col_reg}<19'b0011101010011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011101010011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0011101010011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011101010011101010) && ({row_reg, col_reg}<19'b0011101010011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011101010011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011101010011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011101010011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011101010011101111) && ({row_reg, col_reg}<19'b0011101010100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011101010100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011101010100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0011101010100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0011101010100000100) && ({row_reg, col_reg}<19'b0011101010101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011101010101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0011101010101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011101010110000000) && ({row_reg, col_reg}<19'b0011101010110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011101010110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0011101010110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0011101010110011010) && ({row_reg, col_reg}<19'b0011101100011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011101100011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0011101100011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011101100011101010) && ({row_reg, col_reg}<19'b0011101100011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011101100011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011101100011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011101100011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011101100011101111) && ({row_reg, col_reg}<19'b0011101100100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011101100100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011101100100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0011101100100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0011101100100000100) && ({row_reg, col_reg}<19'b0011101100101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011101100101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0011101100101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011101100110000000) && ({row_reg, col_reg}<19'b0011101100110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011101100110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0011101100110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0011101100110011010) && ({row_reg, col_reg}<19'b0011101110011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011101110011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0011101110011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011101110011101010) && ({row_reg, col_reg}<19'b0011101110011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011101110011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011101110011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011101110011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011101110011101111) && ({row_reg, col_reg}<19'b0011101110100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011101110100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011101110100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0011101110100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0011101110100000100) && ({row_reg, col_reg}<19'b0011101110101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011101110101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0011101110101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011101110110000000) && ({row_reg, col_reg}<19'b0011101110110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011101110110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0011101110110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0011101110110011010) && ({row_reg, col_reg}<19'b0011110000011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011110000011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0011110000011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011110000011101010) && ({row_reg, col_reg}<19'b0011110000011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011110000011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011110000011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011110000011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011110000011101111) && ({row_reg, col_reg}<19'b0011110000100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011110000100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011110000100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0011110000100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0011110000100000100) && ({row_reg, col_reg}<19'b0011110000101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011110000101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0011110000101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011110000110000000) && ({row_reg, col_reg}<19'b0011110000110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011110000110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0011110000110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0011110000110011010) && ({row_reg, col_reg}<19'b0011110010011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011110010011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0011110010011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011110010011101010) && ({row_reg, col_reg}<19'b0011110010011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011110010011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011110010011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011110010011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011110010011101111) && ({row_reg, col_reg}<19'b0011110010100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011110010100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011110010100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0011110010100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0011110010100000100) && ({row_reg, col_reg}<19'b0011110010101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011110010101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0011110010101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011110010110000000) && ({row_reg, col_reg}<19'b0011110010110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011110010110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0011110010110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0011110010110011010) && ({row_reg, col_reg}<19'b0011110100011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011110100011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0011110100011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011110100011101010) && ({row_reg, col_reg}<19'b0011110100011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011110100011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011110100011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011110100011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011110100011101111) && ({row_reg, col_reg}<19'b0011110100100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011110100100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011110100100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0011110100100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0011110100100000100) && ({row_reg, col_reg}<19'b0011110100101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011110100101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0011110100101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011110100110000000) && ({row_reg, col_reg}<19'b0011110100110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011110100110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0011110100110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0011110100110011010) && ({row_reg, col_reg}<19'b0011110110011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011110110011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0011110110011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011110110011101010) && ({row_reg, col_reg}<19'b0011110110011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011110110011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011110110011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011110110011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011110110011101111) && ({row_reg, col_reg}<19'b0011110110100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011110110100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011110110100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0011110110100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0011110110100000100) && ({row_reg, col_reg}<19'b0011110110101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011110110101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0011110110101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011110110110000000) && ({row_reg, col_reg}<19'b0011110110110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011110110110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0011110110110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0011110110110011010) && ({row_reg, col_reg}<19'b0011111000011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011111000011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0011111000011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011111000011101010) && ({row_reg, col_reg}<19'b0011111000011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011111000011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011111000011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011111000011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011111000011101111) && ({row_reg, col_reg}<19'b0011111000100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011111000100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011111000100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0011111000100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0011111000100000100) && ({row_reg, col_reg}<19'b0011111000101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011111000101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0011111000101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011111000110000000) && ({row_reg, col_reg}<19'b0011111000110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011111000110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0011111000110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0011111000110011010) && ({row_reg, col_reg}<19'b0011111010011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011111010011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0011111010011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011111010011101010) && ({row_reg, col_reg}<19'b0011111010011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011111010011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011111010011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011111010011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011111010011101111) && ({row_reg, col_reg}<19'b0011111010100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011111010100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011111010100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0011111010100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0011111010100000100) && ({row_reg, col_reg}<19'b0011111010101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011111010101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0011111010101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011111010110000000) && ({row_reg, col_reg}<19'b0011111010110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011111010110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0011111010110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0011111010110011010) && ({row_reg, col_reg}<19'b0011111100011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011111100011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0011111100011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011111100011101010) && ({row_reg, col_reg}<19'b0011111100011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011111100011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011111100011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011111100011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011111100011101111) && ({row_reg, col_reg}<19'b0011111100100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011111100100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011111100100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0011111100100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0011111100100000100) && ({row_reg, col_reg}<19'b0011111100101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011111100101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0011111100101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011111100110000000) && ({row_reg, col_reg}<19'b0011111100110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011111100110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0011111100110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0011111100110011010) && ({row_reg, col_reg}<19'b0011111110011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011111110011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0011111110011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011111110011101010) && ({row_reg, col_reg}<19'b0011111110011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011111110011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011111110011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011111110011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011111110011101111) && ({row_reg, col_reg}<19'b0011111110100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011111110100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011111110100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0011111110100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0011111110100000100) && ({row_reg, col_reg}<19'b0011111110101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011111110101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0011111110101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011111110110000000) && ({row_reg, col_reg}<19'b0011111110110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011111110110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0011111110110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0011111110110011010) && ({row_reg, col_reg}<19'b0100000000011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100000000011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0100000000011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100000000011101010) && ({row_reg, col_reg}<19'b0100000000011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100000000011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0100000000011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100000000011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100000000011101111) && ({row_reg, col_reg}<19'b0100000000100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100000000100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0100000000100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0100000000100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0100000000100000100) && ({row_reg, col_reg}<19'b0100000000101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100000000101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0100000000101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100000000110000000) && ({row_reg, col_reg}<19'b0100000000110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100000000110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0100000000110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0100000000110011010) && ({row_reg, col_reg}<19'b0100000010011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100000010011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0100000010011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100000010011101010) && ({row_reg, col_reg}<19'b0100000010011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100000010011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0100000010011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100000010011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100000010011101111) && ({row_reg, col_reg}<19'b0100000010100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100000010100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0100000010100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0100000010100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0100000010100000100) && ({row_reg, col_reg}<19'b0100000010101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100000010101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0100000010101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100000010110000000) && ({row_reg, col_reg}<19'b0100000010110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100000010110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0100000010110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0100000010110011010) && ({row_reg, col_reg}<19'b0100000100011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100000100011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0100000100011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100000100011101010) && ({row_reg, col_reg}<19'b0100000100011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100000100011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0100000100011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100000100011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100000100011101111) && ({row_reg, col_reg}<19'b0100000100100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100000100100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0100000100100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0100000100100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0100000100100000100) && ({row_reg, col_reg}<19'b0100000100101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100000100101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0100000100101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100000100110000000) && ({row_reg, col_reg}<19'b0100000100110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100000100110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0100000100110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0100000100110011010) && ({row_reg, col_reg}<19'b0100000110011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100000110011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0100000110011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100000110011101010) && ({row_reg, col_reg}<19'b0100000110011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100000110011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0100000110011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100000110011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100000110011101111) && ({row_reg, col_reg}<19'b0100000110100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100000110100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0100000110100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0100000110100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0100000110100000100) && ({row_reg, col_reg}<19'b0100000110101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100000110101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0100000110101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100000110110000000) && ({row_reg, col_reg}<19'b0100000110110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100000110110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0100000110110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0100000110110011010) && ({row_reg, col_reg}<19'b0100001000011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100001000011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0100001000011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100001000011101010) && ({row_reg, col_reg}<19'b0100001000011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100001000011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0100001000011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100001000011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100001000011101111) && ({row_reg, col_reg}<19'b0100001000100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100001000100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0100001000100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0100001000100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0100001000100000100) && ({row_reg, col_reg}<19'b0100001000101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100001000101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0100001000101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100001000110000000) && ({row_reg, col_reg}<19'b0100001000110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100001000110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0100001000110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0100001000110011010) && ({row_reg, col_reg}<19'b0100001010011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100001010011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0100001010011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100001010011101010) && ({row_reg, col_reg}<19'b0100001010011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100001010011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0100001010011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100001010011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100001010011101111) && ({row_reg, col_reg}<19'b0100001010100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100001010100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0100001010100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0100001010100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0100001010100000100) && ({row_reg, col_reg}<19'b0100001010101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100001010101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0100001010101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100001010110000000) && ({row_reg, col_reg}<19'b0100001010110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100001010110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0100001010110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0100001010110011010) && ({row_reg, col_reg}<19'b0100001100011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100001100011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0100001100011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100001100011101010) && ({row_reg, col_reg}<19'b0100001100011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100001100011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0100001100011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100001100011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100001100011101111) && ({row_reg, col_reg}<19'b0100001100100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100001100100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0100001100100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0100001100100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0100001100100000100) && ({row_reg, col_reg}<19'b0100001100101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100001100101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0100001100101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100001100110000000) && ({row_reg, col_reg}<19'b0100001100110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100001100110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0100001100110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0100001100110011010) && ({row_reg, col_reg}<19'b0100001110011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100001110011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0100001110011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100001110011101010) && ({row_reg, col_reg}<19'b0100001110011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100001110011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0100001110011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100001110011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100001110011101111) && ({row_reg, col_reg}<19'b0100001110100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100001110100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0100001110100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0100001110100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0100001110100000100) && ({row_reg, col_reg}<19'b0100001110101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100001110101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0100001110101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100001110110000000) && ({row_reg, col_reg}<19'b0100001110110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100001110110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0100001110110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0100001110110011010) && ({row_reg, col_reg}<19'b0100010000011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100010000011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0100010000011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100010000011101010) && ({row_reg, col_reg}<19'b0100010000011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100010000011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0100010000011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100010000011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100010000011101111) && ({row_reg, col_reg}<19'b0100010000100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100010000100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0100010000100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0100010000100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0100010000100000100) && ({row_reg, col_reg}<19'b0100010000101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100010000101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0100010000101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100010000110000000) && ({row_reg, col_reg}<19'b0100010000110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100010000110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0100010000110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0100010000110011010) && ({row_reg, col_reg}<19'b0100010010011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100010010011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0100010010011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100010010011101010) && ({row_reg, col_reg}<19'b0100010010011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100010010011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0100010010011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100010010011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100010010011101111) && ({row_reg, col_reg}<19'b0100010010100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100010010100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0100010010100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0100010010100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0100010010100000100) && ({row_reg, col_reg}<19'b0100010010101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100010010101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0100010010101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100010010110000000) && ({row_reg, col_reg}<19'b0100010010110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100010010110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0100010010110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0100010010110011010) && ({row_reg, col_reg}<19'b0100010100011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100010100011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0100010100011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100010100011101010) && ({row_reg, col_reg}<19'b0100010100011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100010100011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0100010100011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100010100011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100010100011101111) && ({row_reg, col_reg}<19'b0100010100100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100010100100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0100010100100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0100010100100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0100010100100000100) && ({row_reg, col_reg}<19'b0100010100101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100010100101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0100010100101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100010100110000000) && ({row_reg, col_reg}<19'b0100010100110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100010100110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0100010100110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0100010100110011010) && ({row_reg, col_reg}<19'b0100010110011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100010110011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0100010110011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100010110011101010) && ({row_reg, col_reg}<19'b0100010110011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100010110011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0100010110011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100010110011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100010110011101111) && ({row_reg, col_reg}<19'b0100010110100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100010110100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0100010110100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0100010110100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0100010110100000100) && ({row_reg, col_reg}<19'b0100010110101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100010110101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0100010110101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100010110110000000) && ({row_reg, col_reg}<19'b0100010110110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100010110110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0100010110110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0100010110110011010) && ({row_reg, col_reg}<19'b0100011000011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100011000011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0100011000011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100011000011101010) && ({row_reg, col_reg}<19'b0100011000011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100011000011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0100011000011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100011000011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100011000011101111) && ({row_reg, col_reg}<19'b0100011000100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100011000100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0100011000100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0100011000100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0100011000100000100) && ({row_reg, col_reg}<19'b0100011000101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100011000101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0100011000101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100011000110000000) && ({row_reg, col_reg}<19'b0100011000110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100011000110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0100011000110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0100011000110011010) && ({row_reg, col_reg}<19'b0100011010011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100011010011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0100011010011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100011010011101010) && ({row_reg, col_reg}<19'b0100011010011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100011010011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0100011010011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100011010011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100011010011101111) && ({row_reg, col_reg}<19'b0100011010100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100011010100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0100011010100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0100011010100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0100011010100000100) && ({row_reg, col_reg}<19'b0100011010101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100011010101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0100011010101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100011010110000000) && ({row_reg, col_reg}<19'b0100011010110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100011010110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0100011010110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0100011010110011010) && ({row_reg, col_reg}<19'b0100011100011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100011100011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0100011100011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100011100011101010) && ({row_reg, col_reg}<19'b0100011100011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100011100011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0100011100011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100011100011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100011100011101111) && ({row_reg, col_reg}<19'b0100011100100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100011100100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0100011100100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0100011100100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0100011100100000100) && ({row_reg, col_reg}<19'b0100011100101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100011100101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0100011100101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100011100110000000) && ({row_reg, col_reg}<19'b0100011100110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100011100110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0100011100110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0100011100110011010) && ({row_reg, col_reg}<19'b0100011110011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100011110011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0100011110011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100011110011101010) && ({row_reg, col_reg}<19'b0100011110011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100011110011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0100011110011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100011110011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100011110011101111) && ({row_reg, col_reg}<19'b0100011110100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100011110100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0100011110100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0100011110100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0100011110100000100) && ({row_reg, col_reg}<19'b0100011110101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100011110101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0100011110101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100011110110000000) && ({row_reg, col_reg}<19'b0100011110110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100011110110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0100011110110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0100011110110011010) && ({row_reg, col_reg}<19'b0100100000011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100100000011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0100100000011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100100000011101010) && ({row_reg, col_reg}<19'b0100100000011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100100000011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0100100000011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100100000011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100100000011101111) && ({row_reg, col_reg}<19'b0100100000100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100100000100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0100100000100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0100100000100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0100100000100000100) && ({row_reg, col_reg}<19'b0100100000101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100100000101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0100100000101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100100000110000000) && ({row_reg, col_reg}<19'b0100100000110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100100000110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0100100000110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0100100000110011010) && ({row_reg, col_reg}<19'b0100100010011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100100010011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0100100010011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100100010011101010) && ({row_reg, col_reg}<19'b0100100010011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100100010011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0100100010011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100100010011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100100010011101111) && ({row_reg, col_reg}<19'b0100100010100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100100010100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0100100010100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0100100010100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0100100010100000100) && ({row_reg, col_reg}<19'b0100100010101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100100010101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0100100010101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100100010110000000) && ({row_reg, col_reg}<19'b0100100010110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100100010110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0100100010110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0100100010110011010) && ({row_reg, col_reg}<19'b0100100100011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100100100011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0100100100011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100100100011101010) && ({row_reg, col_reg}<19'b0100100100011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100100100011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0100100100011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100100100011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100100100011101111) && ({row_reg, col_reg}<19'b0100100100100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100100100100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0100100100100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0100100100100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0100100100100000100) && ({row_reg, col_reg}<19'b0100100100101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100100100101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0100100100101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100100100110000000) && ({row_reg, col_reg}<19'b0100100100110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100100100110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0100100100110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0100100100110011010) && ({row_reg, col_reg}<19'b0100100110011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100100110011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0100100110011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100100110011101010) && ({row_reg, col_reg}<19'b0100100110011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100100110011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0100100110011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100100110011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100100110011101111) && ({row_reg, col_reg}<19'b0100100110100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100100110100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0100100110100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0100100110100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0100100110100000100) && ({row_reg, col_reg}<19'b0100100110101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100100110101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0100100110101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100100110110000000) && ({row_reg, col_reg}<19'b0100100110110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100100110110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0100100110110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0100100110110011010) && ({row_reg, col_reg}<19'b0100101000011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100101000011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0100101000011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100101000011101010) && ({row_reg, col_reg}<19'b0100101000011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100101000011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0100101000011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100101000011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100101000011101111) && ({row_reg, col_reg}<19'b0100101000100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100101000100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0100101000100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0100101000100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0100101000100000100) && ({row_reg, col_reg}<19'b0100101000101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100101000101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0100101000101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100101000110000000) && ({row_reg, col_reg}<19'b0100101000110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100101000110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0100101000110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0100101000110011010) && ({row_reg, col_reg}<19'b0100101010011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100101010011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0100101010011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100101010011101010) && ({row_reg, col_reg}<19'b0100101010011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100101010011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0100101010011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100101010011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100101010011101111) && ({row_reg, col_reg}<19'b0100101010100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100101010100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0100101010100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0100101010100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0100101010100000100) && ({row_reg, col_reg}<19'b0100101010101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100101010101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0100101010101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100101010110000000) && ({row_reg, col_reg}<19'b0100101010110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100101010110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0100101010110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0100101010110011010) && ({row_reg, col_reg}<19'b0100101100011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100101100011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0100101100011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100101100011101010) && ({row_reg, col_reg}<19'b0100101100011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100101100011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0100101100011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100101100011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100101100011101111) && ({row_reg, col_reg}<19'b0100101100100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100101100100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0100101100100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0100101100100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0100101100100000100) && ({row_reg, col_reg}<19'b0100101100101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100101100101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0100101100101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100101100110000000) && ({row_reg, col_reg}<19'b0100101100110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100101100110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0100101100110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0100101100110011010) && ({row_reg, col_reg}<19'b0100101110011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100101110011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0100101110011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100101110011101010) && ({row_reg, col_reg}<19'b0100101110011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100101110011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0100101110011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100101110011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100101110011101111) && ({row_reg, col_reg}<19'b0100101110100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100101110100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0100101110100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0100101110100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0100101110100000100) && ({row_reg, col_reg}<19'b0100101110101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100101110101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0100101110101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100101110110000000) && ({row_reg, col_reg}<19'b0100101110110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100101110110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0100101110110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0100101110110011010) && ({row_reg, col_reg}<19'b0100110000011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100110000011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0100110000011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100110000011101010) && ({row_reg, col_reg}<19'b0100110000011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100110000011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0100110000011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100110000011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100110000011101111) && ({row_reg, col_reg}<19'b0100110000100000000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0100110000100000000) && ({row_reg, col_reg}<19'b0100110000100000010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0100110000100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0100110000100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0100110000100000100) && ({row_reg, col_reg}<19'b0100110000101111101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100110000101111101)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0100110000101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0100110000101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100110000110000000) && ({row_reg, col_reg}<19'b0100110000110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100110000110011000)) color_data = 12'b101010101010;

		if(({row_reg, col_reg}>=19'b0100110000110011001) && ({row_reg, col_reg}<19'b0100110010011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100110010011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0100110010011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100110010011101010) && ({row_reg, col_reg}<19'b0100110010011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100110010011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0100110010011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100110010011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100110010011101111) && ({row_reg, col_reg}<19'b0100110010100000010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100110010100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0100110010100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0100110010100000100) && ({row_reg, col_reg}<19'b0100110010101111101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100110010101111101)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0100110010101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0100110010101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100110010110000000) && ({row_reg, col_reg}<19'b0100110010110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100110010110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0100110010110011001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=19'b0100110010110011010) && ({row_reg, col_reg}<19'b0100110011000101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100110011000101000)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0100110011000101001) && ({row_reg, col_reg}<19'b0100110100001011100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100110100001011100)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=19'b0100110100001011101) && ({row_reg, col_reg}<19'b0100110100001100000)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0100110100001100000) && ({row_reg, col_reg}<19'b0100110100011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0100110100011101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0100110100011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100110100011101010) && ({row_reg, col_reg}<19'b0100110100011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100110100011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0100110100011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100110100011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100110100011101111) && ({row_reg, col_reg}<19'b0100110100100000000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0100110100100000000) && ({row_reg, col_reg}<19'b0100110100100000010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0100110100100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0100110100100000011)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=19'b0100110100100000100) && ({row_reg, col_reg}<19'b0100110100101111100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0100110100101111100)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0100110100101111101)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0100110100101111110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0100110100101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100110100110000000) && ({row_reg, col_reg}<19'b0100110100110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100110100110011000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=19'b0100110100110011001) && ({row_reg, col_reg}<19'b0100110101000100011)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=19'b0100110101000100011) && ({row_reg, col_reg}<19'b0100110101000100101)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0100110101000100101)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0100110101000100110) && ({row_reg, col_reg}<19'b0100110110001011001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100110110001011001)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0100110110001011010) && ({row_reg, col_reg}<19'b0100110110001011100)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0100110110001011100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=19'b0100110110001011101) && ({row_reg, col_reg}<19'b0100110110001011111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=19'b0100110110001011111) && ({row_reg, col_reg}<19'b0100110110011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0100110110011101001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100110110011101010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0100110110011101011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100110110011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100110110011101101) && ({row_reg, col_reg}<19'b0100110110011101111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100110110011101111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100110110011110000) && ({row_reg, col_reg}<19'b0100110110100000011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0100110110100000011) && ({row_reg, col_reg}<19'b0100110110101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100110110101111111) && ({row_reg, col_reg}<19'b0100110110110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100110110110011000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0100110110110011001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=19'b0100110110110011010) && ({row_reg, col_reg}<19'b0100110110110011101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100110110110011101) && ({row_reg, col_reg}<19'b0100110110110011111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=19'b0100110110110011111) && ({row_reg, col_reg}<19'b0100110111000100011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100110111000100011) && ({row_reg, col_reg}<19'b0100110111000100101)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0100110111000100101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0100110111000100110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0100110111000100111)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0100110111000101000)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0100110111000101001) && ({row_reg, col_reg}<19'b0100111000001010111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100111000001010111)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0100111000001011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0100111000001011001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=19'b0100111000001011010) && ({row_reg, col_reg}<19'b0100111000001011100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100111000001011100) && ({row_reg, col_reg}<19'b0100111000001011110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0100111000001011110) && ({row_reg, col_reg}<19'b0100111000001100000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100111000001100000) && ({row_reg, col_reg}<19'b0100111000011101010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100111000011101010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100111000011101011) && ({row_reg, col_reg}<19'b0100111000100000000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0100111000100000000) && ({row_reg, col_reg}<19'b0100111000100000010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0100111000100000010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100111000100000011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0100111000100000100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0100111000100000101) && ({row_reg, col_reg}<19'b0100111000100001000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100111000100001000) && ({row_reg, col_reg}<19'b0100111000101111000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0100111000101111000) && ({row_reg, col_reg}<19'b0100111000101111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0100111000101111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0100111000101111101) && ({row_reg, col_reg}<19'b0100111000101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100111000101111111) && ({row_reg, col_reg}<19'b0100111000110011101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100111000110011101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100111000110011110) && ({row_reg, col_reg}<19'b0100111001000100000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100111001000100000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100111001000100001) && ({row_reg, col_reg}<19'b0100111001000100011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100111001000100011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100111001000100100) && ({row_reg, col_reg}<19'b0100111001000100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0100111001000100110) && ({row_reg, col_reg}<19'b0100111001000101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0100111001000101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0100111001000101001)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=19'b0100111001000101010) && ({row_reg, col_reg}<19'b0100111010001010101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100111010001010101)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0100111010001010110)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0100111010001010111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0100111010001011000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100111010001011001) && ({row_reg, col_reg}<19'b0100111010001011011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0100111010001011011) && ({row_reg, col_reg}<19'b0100111010001011111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100111010001011111) && ({row_reg, col_reg}<19'b0100111010011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0100111010011101101) && ({row_reg, col_reg}<19'b0100111010011101111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100111010011101111) && ({row_reg, col_reg}<19'b0100111010100000000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0100111010100000000) && ({row_reg, col_reg}<19'b0100111010100000010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100111010100000010) && ({row_reg, col_reg}<19'b0100111010101111011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100111010101111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0100111010101111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0100111010101111101) && ({row_reg, col_reg}<19'b0100111010101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100111010101111111) && ({row_reg, col_reg}<19'b0100111010110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0100111010110011000) && ({row_reg, col_reg}<19'b0100111010110011100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100111010110011100) && ({row_reg, col_reg}<19'b0100111010110011111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100111010110011111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100111010110100000) && ({row_reg, col_reg}<19'b0100111011000100100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100111011000100100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100111011000100101) && ({row_reg, col_reg}<19'b0100111011000101001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100111011000101001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0100111011000101010)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0100111011000101011)) color_data = 12'b110111011101;

		if(({row_reg, col_reg}>=19'b0100111011000101100) && ({row_reg, col_reg}<19'b0100111100001010100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100111100001010100)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0100111100001010101)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0100111100001010110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=19'b0100111100001010111) && ({row_reg, col_reg}<19'b0100111100001011110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100111100001011110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100111100001011111) && ({row_reg, col_reg}<19'b0100111100011101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100111100011101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100111100011101001) && ({row_reg, col_reg}<19'b0100111100011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0100111100011101101) && ({row_reg, col_reg}<19'b0100111100011101111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100111100011101111) && ({row_reg, col_reg}<19'b0100111100100000010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100111100100000010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0100111100100000011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0100111100100000100) && ({row_reg, col_reg}<19'b0100111100100001000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100111100100001000) && ({row_reg, col_reg}<19'b0100111100101111000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0100111100101111000) && ({row_reg, col_reg}<19'b0100111100101111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0100111100101111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100111100101111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100111100101111100) && ({row_reg, col_reg}<19'b0100111100110011010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100111100110011010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100111100110011011) && ({row_reg, col_reg}<19'b0100111100110011111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100111100110011111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100111100110100000) && ({row_reg, col_reg}<19'b0100111101000100000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0100111101000100000) && ({row_reg, col_reg}<19'b0100111101000100011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100111101000100011) && ({row_reg, col_reg}<19'b0100111101000101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100111101000101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0100111101000101001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100111101000101010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0100111101000101011)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0100111101000101100)) color_data = 12'b110111011101;

		if(({row_reg, col_reg}>=19'b0100111101000101101) && ({row_reg, col_reg}<19'b0100111110001010100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100111110001010100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0100111110001010101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0100111110001010110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100111110001010111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0100111110001011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0100111110001011001) && ({row_reg, col_reg}<19'b0100111110001011101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100111110001011101) && ({row_reg, col_reg}<19'b0100111110011101001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100111110011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0100111110011101010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100111110011101011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100111110011101100) && ({row_reg, col_reg}<19'b0100111110100000000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100111110100000000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100111110100000001) && ({row_reg, col_reg}<19'b0100111110100000101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100111110100000101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100111110100000110) && ({row_reg, col_reg}<19'b0100111110101111011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100111110101111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100111110101111100) && ({row_reg, col_reg}<19'b0100111110101111111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100111110101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100111110110000000) && ({row_reg, col_reg}<19'b0100111110110011100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0100111110110011100) && ({row_reg, col_reg}<19'b0100111110110011110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100111110110011110) && ({row_reg, col_reg}<19'b0100111111000100010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0100111111000100010) && ({row_reg, col_reg}<19'b0100111111000100100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100111111000100100) && ({row_reg, col_reg}<19'b0100111111000100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0100111111000100110) && ({row_reg, col_reg}<19'b0100111111000101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0100111111000101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100111111000101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0100111111000101010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100111111000101011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0100111111000101100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0100111111000101101)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0100111111000101110) && ({row_reg, col_reg}<19'b0101000000001010011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101000000001010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0101000000001010100)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=19'b0101000000001010101) && ({row_reg, col_reg}<19'b0101000001000101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0101000001000101000) && ({row_reg, col_reg}<19'b0101000001000101010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101000001000101010) && ({row_reg, col_reg}<19'b0101000001000101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101000001000101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101000001000101101)) color_data = 12'b101110111011;

		if(({row_reg, col_reg}>=19'b0101000001000101110) && ({row_reg, col_reg}<19'b0101000010001010010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101000010001010010)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0101000010001010011)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0101000010001010100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101000010001010101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101000010001010110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101000010001010111) && ({row_reg, col_reg}<19'b0101000011000101001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0101000011000101001) && ({row_reg, col_reg}<19'b0101000011000101011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101000011000101011) && ({row_reg, col_reg}<19'b0101000011000101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101000011000101101)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0101000011000101110)) color_data = 12'b110111011101;

		if(({row_reg, col_reg}>=19'b0101000011000101111) && ({row_reg, col_reg}<19'b0101000100001010010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101000100001010010)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0101000100001010011)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=19'b0101000100001010100) && ({row_reg, col_reg}<19'b0101000100001010110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101000100001010110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101000100001010111) && ({row_reg, col_reg}<19'b0101000101000101001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0101000101000101001) && ({row_reg, col_reg}<19'b0101000101000101011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101000101000101011) && ({row_reg, col_reg}<19'b0101000101000101110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101000101000101110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0101000101000101111)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0101000101000110000) && ({row_reg, col_reg}<19'b0101000110001010001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101000110001010001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0101000110001010010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0101000110001010011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101000110001010100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101000110001010101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101000110001010110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101000110001010111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101000110001011000) && ({row_reg, col_reg}<19'b0101000111000101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101000111000101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101000111000101001) && ({row_reg, col_reg}<19'b0101000111000101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101000111000101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101000111000101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101000111000101110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0101000111000101111)) color_data = 12'b110111011101;

		if(({row_reg, col_reg}>=19'b0101000111000110000) && ({row_reg, col_reg}<19'b0101001000001010001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101001000001010001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0101001000001010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0101001000001010011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101001000001010100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101001000001010101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101001000001010110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101001000001010111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101001000001011000) && ({row_reg, col_reg}<19'b0101001001000101010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101001001000101010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101001001000101011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101001001000101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101001001000101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101001001000101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101001001000101111)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=19'b0101001001000110000) && ({row_reg, col_reg}<19'b0101001010001010001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101001010001010001)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0101001010001010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=19'b0101001010001010011) && ({row_reg, col_reg}<19'b0101001010001010101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101001010001010101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101001010001010110) && ({row_reg, col_reg}<19'b0101001011000101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101001011000101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101001011000101001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101001011000101010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101001011000101011) && ({row_reg, col_reg}<19'b0101001011000101110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101001011000101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101001011000101111)) color_data = 12'b101010101010;

		if(({row_reg, col_reg}>=19'b0101001011000110000) && ({row_reg, col_reg}<19'b0101001100001010001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101001100001010001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0101001100001010010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101001100001010011) && ({row_reg, col_reg}<19'b0101001100001010101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101001100001010101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101001100001010110) && ({row_reg, col_reg}<19'b0101001101000101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101001101000101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101001101000101001) && ({row_reg, col_reg}<19'b0101001101000101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0101001101000101101) && ({row_reg, col_reg}<19'b0101001101000101111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101001101000101111)) color_data = 12'b100110011001;

		if(({row_reg, col_reg}>=19'b0101001101000110000) && ({row_reg, col_reg}<19'b0101001110001010001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101001110001010001)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=19'b0101001110001010010) && ({row_reg, col_reg}<19'b0101001110001010100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101001110001010100) && ({row_reg, col_reg}<19'b0101001110001010111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101001110001010111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101001110001011000) && ({row_reg, col_reg}<19'b0101001111000101010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0101001111000101010) && ({row_reg, col_reg}<19'b0101001111000101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101001111000101100) && ({row_reg, col_reg}<19'b0101001111000101111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101001111000101111)) color_data = 12'b100010001000;

		if(({row_reg, col_reg}>=19'b0101001111000110000) && ({row_reg, col_reg}<19'b0101010000001010001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101010000001010001)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0101010000001010010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101010000001010011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101010000001010100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101010000001010101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101010000001010110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101010000001010111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101010000001011000) && ({row_reg, col_reg}<19'b0101010001000101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101010001000101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101010001000101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101010001000101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101010001000101111)) color_data = 12'b100110011001;

		if(({row_reg, col_reg}>=19'b0101010001000110000) && ({row_reg, col_reg}<19'b0101010010001010001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101010010001010001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=19'b0101010010001010010) && ({row_reg, col_reg}<19'b0101010010001010100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101010010001010100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101010010001010101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101010010001010110) && ({row_reg, col_reg}<19'b0101010011000101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0101010011000101000) && ({row_reg, col_reg}<19'b0101010011000101011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101010011000101011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101010011000101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101010011000101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101010011000101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101010011000101111)) color_data = 12'b101010101010;

		if(({row_reg, col_reg}>=19'b0101010011000110000) && ({row_reg, col_reg}<19'b0101010100001010001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101010100001010001)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0101010100001010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0101010100001010011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0101010100001010100) && ({row_reg, col_reg}<19'b0101010100001010110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101010100001010110) && ({row_reg, col_reg}<19'b0101010101000101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101010101000101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101010101000101001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101010101000101010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101010101000101011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101010101000101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101010101000101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101010101000101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101010101000101111)) color_data = 12'b101110111011;

		if(({row_reg, col_reg}>=19'b0101010101000110000) && ({row_reg, col_reg}<19'b0101010110001010001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101010110001010001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0101010110001010010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0101010110001010011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0101010110001010100) && ({row_reg, col_reg}<19'b0101010110001010110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101010110001010110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101010110001010111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101010110001011000) && ({row_reg, col_reg}<19'b0101010111000101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101010111000101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101010111000101001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101010111000101010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101010111000101011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101010111000101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101010111000101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101010111000101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101010111000101111)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=19'b0101010111000110000) && ({row_reg, col_reg}<19'b0101011000001010010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101011000001010010)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0101011000001010011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101011000001010100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101011000001010101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101011000001010110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101011000001010111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101011000001011000) && ({row_reg, col_reg}<19'b0101011001000101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101011001000101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101011001000101001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0101011001000101010) && ({row_reg, col_reg}<19'b0101011001000101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101011001000101100) && ({row_reg, col_reg}<19'b0101011001000101110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101011001000101110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0101011001000101111)) color_data = 12'b110111011101;

		if(({row_reg, col_reg}>=19'b0101011001000110000) && ({row_reg, col_reg}<19'b0101011010001010010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101011010001010010)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0101011010001010011)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=19'b0101011010001010100) && ({row_reg, col_reg}<19'b0101011011000101010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0101011011000101010) && ({row_reg, col_reg}<19'b0101011011000101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101011011000101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101011011000101101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101011011000101110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0101011011000101111)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0101011011000110000) && ({row_reg, col_reg}<19'b0101011100001010010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101011100001010010)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0101011100001010011)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0101011100001010100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101011100001010101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101011100001010110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101011100001010111) && ({row_reg, col_reg}<19'b0101011101000101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101011101000101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101011101000101101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0101011101000101110)) color_data = 12'b110111011101;

		if(({row_reg, col_reg}>=19'b0101011101000101111) && ({row_reg, col_reg}<19'b0101011110001010011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101011110001010011)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0101011110001010100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=19'b0101011110001010101) && ({row_reg, col_reg}<19'b0101011110001010111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101011110001010111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101011110001011000) && ({row_reg, col_reg}<19'b0101011111000101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0101011111000101000) && ({row_reg, col_reg}<19'b0101011111000101010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101011111000101010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0101011111000101011) && ({row_reg, col_reg}<19'b0101011111000101101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101011111000101101)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=19'b0101011111000101110) && ({row_reg, col_reg}<19'b0101100000001010100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101100000001010100)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0101100000001010101)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=19'b0101100000001010110) && ({row_reg, col_reg}<19'b0101100000001011101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0101100000001011101) && ({row_reg, col_reg}<19'b0101100000001011111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101100000001011111) && ({row_reg, col_reg}<19'b0101100000011101010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101100000011101010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101100000011101011) && ({row_reg, col_reg}<19'b0101100000011101111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101100000011101111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101100000011110000) && ({row_reg, col_reg}<19'b0101100000100000000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101100000100000000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101100000100000001) && ({row_reg, col_reg}<19'b0101100000100000100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101100000100000100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101100000100000101) && ({row_reg, col_reg}<19'b0101100000100000111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101100000100000111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101100000100001000) && ({row_reg, col_reg}<19'b0101100000101111000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101100000101111000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101100000101111001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101100000101111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101100000101111011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101100000101111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101100000101111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101100000101111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101100000101111111) && ({row_reg, col_reg}<19'b0101100000110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0101100000110011000) && ({row_reg, col_reg}<19'b0101100000110011010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101100000110011010) && ({row_reg, col_reg}<19'b0101100000110011101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101100000110011101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101100000110011110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101100000110011111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101100000110100000) && ({row_reg, col_reg}<19'b0101100001000100000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0101100001000100000) && ({row_reg, col_reg}<19'b0101100001000100010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101100001000100010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0101100001000100011) && ({row_reg, col_reg}<19'b0101100001000100110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101100001000100110) && ({row_reg, col_reg}<19'b0101100001000101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101100001000101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101100001000101001) && ({row_reg, col_reg}<19'b0101100001000101011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101100001000101011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101100001000101100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0101100001000101101)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0101100001000101110) && ({row_reg, col_reg}<19'b0101100010001010100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101100010001010100)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0101100010001010101)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0101100010001010110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0101100010001010111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101100010001011000) && ({row_reg, col_reg}<19'b0101100010001011010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0101100010001011010) && ({row_reg, col_reg}<19'b0101100010001011100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101100010001011100) && ({row_reg, col_reg}<19'b0101100010011101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101100010011101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101100010011101001) && ({row_reg, col_reg}<19'b0101100010100000010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101100010100000010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101100010100000011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0101100010100000100) && ({row_reg, col_reg}<19'b0101100010100000110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101100010100000110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101100010100000111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101100010100001000) && ({row_reg, col_reg}<19'b0101100010101111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101100010101111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101100010101111011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0101100010101111100) && ({row_reg, col_reg}<19'b0101100010101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101100010101111111) && ({row_reg, col_reg}<19'b0101100010110011001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0101100010110011001) && ({row_reg, col_reg}<19'b0101100010110011011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101100010110011011) && ({row_reg, col_reg}<19'b0101100010110011101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101100010110011101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101100010110011110) && ({row_reg, col_reg}<19'b0101100011000100000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101100011000100000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101100011000100001) && ({row_reg, col_reg}<19'b0101100011000100101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0101100011000100101) && ({row_reg, col_reg}<19'b0101100011000101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101100011000101000) && ({row_reg, col_reg}<19'b0101100011000101010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101100011000101010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0101100011000101011)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0101100011000101100)) color_data = 12'b110111011101;

		if(({row_reg, col_reg}>=19'b0101100011000101101) && ({row_reg, col_reg}<19'b0101100100001010110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101100100001010110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0101100100001010111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=19'b0101100100001011000) && ({row_reg, col_reg}<19'b0101100100001011010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101100100001011010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0101100100001011011) && ({row_reg, col_reg}<19'b0101100100011101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101100100011101000) && ({row_reg, col_reg}<19'b0101100100011101010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101100100011101010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101100100011101011) && ({row_reg, col_reg}<19'b0101100100011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101100100011101101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101100100011101110) && ({row_reg, col_reg}<19'b0101100100100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0101100100100000001) && ({row_reg, col_reg}<19'b0101100100100000011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101100100100000011) && ({row_reg, col_reg}<19'b0101100100100001000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0101100100100001000) && ({row_reg, col_reg}<19'b0101100100101111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101100100101111001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101100100101111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101100100101111011) && ({row_reg, col_reg}<19'b0101100100110011001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0101100100110011001) && ({row_reg, col_reg}<19'b0101100100110011100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101100100110011100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0101100100110011101) && ({row_reg, col_reg}<19'b0101100100110011111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101100100110011111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0101100100110100000) && ({row_reg, col_reg}<19'b0101100101000100000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101100101000100000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0101100101000100001) && ({row_reg, col_reg}<19'b0101100101000100101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101100101000100101) && ({row_reg, col_reg}<19'b0101100101000101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101100101000101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101100101000101001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0101100101000101010)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0101100101000101011)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0101100101000101100) && ({row_reg, col_reg}<19'b0101100110001010111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101100110001010111)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0101100110001011000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0101100110001011001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=19'b0101100110001011010) && ({row_reg, col_reg}<19'b0101100110001011100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101100110001011100) && ({row_reg, col_reg}<19'b0101100110011101010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101100110011101010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101100110011101011) && ({row_reg, col_reg}<19'b0101100110011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101100110011101101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101100110011101110) && ({row_reg, col_reg}<19'b0101100110100000101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0101100110100000101) && ({row_reg, col_reg}<19'b0101100110100001000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101100110100001000) && ({row_reg, col_reg}<19'b0101100110101111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101100110101111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101100110101111011) && ({row_reg, col_reg}<19'b0101100110101111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0101100110101111101) && ({row_reg, col_reg}<19'b0101100110110000000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101100110110000000) && ({row_reg, col_reg}<19'b0101100110110011001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101100110110011001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101100110110011010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101100110110011011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101100110110011100) && ({row_reg, col_reg}<19'b0101100111000100101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0101100111000100101) && ({row_reg, col_reg}<19'b0101100111000100111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101100111000100111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0101100111000101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0101100111000101001)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0101100111000101010)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0101100111000101011) && ({row_reg, col_reg}<19'b0101101000001011001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101101000001011001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0101101000001011010)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=19'b0101101000001011011) && ({row_reg, col_reg}<19'b0101101000001011101)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0101101000001011101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=19'b0101101000001011110) && ({row_reg, col_reg}<19'b0101101000011101001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=19'b0101101000011101001) && ({row_reg, col_reg}<19'b0101101000011101011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101101000011101011) && ({row_reg, col_reg}<19'b0101101000011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101101000011101101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101101000011101110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101101000011101111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101101000011110000) && ({row_reg, col_reg}<19'b0101101000100000000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0101101000100000000) && ({row_reg, col_reg}<19'b0101101000100000011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101101000100000011) && ({row_reg, col_reg}<19'b0101101000101111110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0101101000101111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101101000101111111) && ({row_reg, col_reg}<19'b0101101000110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101101000110011000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101101000110011001) && ({row_reg, col_reg}<19'b0101101001000100100)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0101101001000100100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0101101001000100101)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0101101001000100110)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0101101001000100111)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0101101001000101000)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0101101001000101001) && ({row_reg, col_reg}<19'b0101101010001011101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101101010001011101)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=19'b0101101010001011110) && ({row_reg, col_reg}<19'b0101101010011101000)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0101101010011101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0101101010011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101101010011101010) && ({row_reg, col_reg}<19'b0101101010011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101101010011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101101010011101101) && ({row_reg, col_reg}<19'b0101101010011101111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101101010011101111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101101010011110000) && ({row_reg, col_reg}<19'b0101101010100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101101010100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101101010100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0101101010100000011)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=19'b0101101010100000100) && ({row_reg, col_reg}<19'b0101101010100000111)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0101101010100000111)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=19'b0101101010100001000) && ({row_reg, col_reg}<19'b0101101010101111000)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0101101010101111000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=19'b0101101010101111001) && ({row_reg, col_reg}<19'b0101101010101111110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0101101010101111110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0101101010101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101101010110000000) && ({row_reg, col_reg}<19'b0101101010110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101101010110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=19'b0101101010110011001) && ({row_reg, col_reg}<19'b0101101011000100011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0101101011000100011) && ({row_reg, col_reg}<19'b0101101011000100101)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0101101011000100101) && ({row_reg, col_reg}<19'b0101101100011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101101100011101000)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0101101100011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101101100011101010) && ({row_reg, col_reg}<19'b0101101100011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101101100011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101101100011101101) && ({row_reg, col_reg}<19'b0101101100011101111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101101100011101111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101101100011110000) && ({row_reg, col_reg}<19'b0101101100100000010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101101100100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0101101100100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0101101100100000100) && ({row_reg, col_reg}<19'b0101101100101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101101100101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0101101100101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101101100110000000) && ({row_reg, col_reg}<19'b0101101100110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101101100110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0101101100110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0101101100110011010) && ({row_reg, col_reg}<19'b0101101110011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101101110011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=19'b0101101110011101001) && ({row_reg, col_reg}<19'b0101101110011101011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101101110011101011) && ({row_reg, col_reg}<19'b0101101110011101110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101101110011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101101110011101111) && ({row_reg, col_reg}<19'b0101101110100000000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101101110100000000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101101110100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101101110100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0101101110100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0101101110100000100) && ({row_reg, col_reg}<19'b0101101110101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101101110101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0101101110101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101101110110000000) && ({row_reg, col_reg}<19'b0101101110110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101101110110011000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0101101110110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0101101110110011010) && ({row_reg, col_reg}<19'b0101110000011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101110000011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0101110000011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101110000011101010) && ({row_reg, col_reg}<19'b0101110000011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101110000011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101110000011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101110000011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101110000011101111) && ({row_reg, col_reg}<19'b0101110000100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101110000100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101110000100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0101110000100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0101110000100000100) && ({row_reg, col_reg}<19'b0101110000101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101110000101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0101110000101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101110000110000000) && ({row_reg, col_reg}<19'b0101110000110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101110000110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0101110000110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0101110000110011010) && ({row_reg, col_reg}<19'b0101110010011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101110010011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0101110010011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101110010011101010) && ({row_reg, col_reg}<19'b0101110010011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101110010011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101110010011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101110010011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101110010011101111) && ({row_reg, col_reg}<19'b0101110010100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101110010100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101110010100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0101110010100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0101110010100000100) && ({row_reg, col_reg}<19'b0101110010101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101110010101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0101110010101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101110010110000000) && ({row_reg, col_reg}<19'b0101110010110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101110010110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0101110010110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0101110010110011010) && ({row_reg, col_reg}<19'b0101110100011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101110100011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0101110100011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101110100011101010) && ({row_reg, col_reg}<19'b0101110100011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101110100011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101110100011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101110100011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101110100011101111) && ({row_reg, col_reg}<19'b0101110100100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101110100100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101110100100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0101110100100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0101110100100000100) && ({row_reg, col_reg}<19'b0101110100101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101110100101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0101110100101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101110100110000000) && ({row_reg, col_reg}<19'b0101110100110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101110100110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0101110100110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0101110100110011010) && ({row_reg, col_reg}<19'b0101110110011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101110110011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0101110110011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101110110011101010) && ({row_reg, col_reg}<19'b0101110110011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101110110011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101110110011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101110110011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101110110011101111) && ({row_reg, col_reg}<19'b0101110110100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101110110100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101110110100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0101110110100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0101110110100000100) && ({row_reg, col_reg}<19'b0101110110101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101110110101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0101110110101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101110110110000000) && ({row_reg, col_reg}<19'b0101110110110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101110110110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0101110110110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0101110110110011010) && ({row_reg, col_reg}<19'b0101111000011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101111000011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0101111000011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101111000011101010) && ({row_reg, col_reg}<19'b0101111000011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101111000011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101111000011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101111000011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101111000011101111) && ({row_reg, col_reg}<19'b0101111000100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101111000100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101111000100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0101111000100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0101111000100000100) && ({row_reg, col_reg}<19'b0101111000101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101111000101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0101111000101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101111000110000000) && ({row_reg, col_reg}<19'b0101111000110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101111000110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0101111000110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0101111000110011010) && ({row_reg, col_reg}<19'b0101111010011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101111010011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0101111010011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101111010011101010) && ({row_reg, col_reg}<19'b0101111010011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101111010011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101111010011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101111010011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101111010011101111) && ({row_reg, col_reg}<19'b0101111010100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101111010100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101111010100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0101111010100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0101111010100000100) && ({row_reg, col_reg}<19'b0101111010101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101111010101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0101111010101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101111010110000000) && ({row_reg, col_reg}<19'b0101111010110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101111010110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0101111010110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0101111010110011010) && ({row_reg, col_reg}<19'b0101111100011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101111100011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0101111100011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101111100011101010) && ({row_reg, col_reg}<19'b0101111100011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101111100011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101111100011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101111100011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101111100011101111) && ({row_reg, col_reg}<19'b0101111100100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101111100100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101111100100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0101111100100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0101111100100000100) && ({row_reg, col_reg}<19'b0101111100101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101111100101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0101111100101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101111100110000000) && ({row_reg, col_reg}<19'b0101111100110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101111100110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0101111100110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0101111100110011010) && ({row_reg, col_reg}<19'b0101111110011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101111110011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0101111110011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101111110011101010) && ({row_reg, col_reg}<19'b0101111110011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101111110011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101111110011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101111110011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101111110011101111) && ({row_reg, col_reg}<19'b0101111110100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101111110100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101111110100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0101111110100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0101111110100000100) && ({row_reg, col_reg}<19'b0101111110101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101111110101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0101111110101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101111110110000000) && ({row_reg, col_reg}<19'b0101111110110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101111110110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0101111110110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0101111110110011010) && ({row_reg, col_reg}<19'b0110000000011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0110000000011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0110000000011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0110000000011101010) && ({row_reg, col_reg}<19'b0110000000011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110000000011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0110000000011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110000000011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0110000000011101111) && ({row_reg, col_reg}<19'b0110000000100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110000000100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0110000000100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0110000000100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0110000000100000100) && ({row_reg, col_reg}<19'b0110000000101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0110000000101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0110000000101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0110000000110000000) && ({row_reg, col_reg}<19'b0110000000110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110000000110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0110000000110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0110000000110011010) && ({row_reg, col_reg}<19'b0110000010011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0110000010011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0110000010011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0110000010011101010) && ({row_reg, col_reg}<19'b0110000010011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110000010011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0110000010011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110000010011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0110000010011101111) && ({row_reg, col_reg}<19'b0110000010100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110000010100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0110000010100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0110000010100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0110000010100000100) && ({row_reg, col_reg}<19'b0110000010101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0110000010101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0110000010101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0110000010110000000) && ({row_reg, col_reg}<19'b0110000010110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110000010110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0110000010110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0110000010110011010) && ({row_reg, col_reg}<19'b0110000100011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0110000100011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0110000100011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0110000100011101010) && ({row_reg, col_reg}<19'b0110000100011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110000100011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0110000100011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110000100011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0110000100011101111) && ({row_reg, col_reg}<19'b0110000100100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110000100100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0110000100100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0110000100100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0110000100100000100) && ({row_reg, col_reg}<19'b0110000100101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0110000100101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0110000100101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0110000100110000000) && ({row_reg, col_reg}<19'b0110000100110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110000100110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0110000100110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0110000100110011010) && ({row_reg, col_reg}<19'b0110000110011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0110000110011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0110000110011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0110000110011101010) && ({row_reg, col_reg}<19'b0110000110011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110000110011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0110000110011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110000110011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0110000110011101111) && ({row_reg, col_reg}<19'b0110000110100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110000110100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0110000110100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0110000110100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0110000110100000100) && ({row_reg, col_reg}<19'b0110000110101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0110000110101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0110000110101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0110000110110000000) && ({row_reg, col_reg}<19'b0110000110110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110000110110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0110000110110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0110000110110011010) && ({row_reg, col_reg}<19'b0110001000011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0110001000011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0110001000011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0110001000011101010) && ({row_reg, col_reg}<19'b0110001000011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110001000011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0110001000011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110001000011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0110001000011101111) && ({row_reg, col_reg}<19'b0110001000100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110001000100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0110001000100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0110001000100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0110001000100000100) && ({row_reg, col_reg}<19'b0110001000101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0110001000101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0110001000101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0110001000110000000) && ({row_reg, col_reg}<19'b0110001000110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110001000110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0110001000110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0110001000110011010) && ({row_reg, col_reg}<19'b0110001010011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0110001010011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0110001010011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0110001010011101010) && ({row_reg, col_reg}<19'b0110001010011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110001010011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0110001010011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110001010011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0110001010011101111) && ({row_reg, col_reg}<19'b0110001010100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110001010100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0110001010100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0110001010100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0110001010100000100) && ({row_reg, col_reg}<19'b0110001010101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0110001010101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0110001010101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0110001010110000000) && ({row_reg, col_reg}<19'b0110001010110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110001010110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0110001010110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0110001010110011010) && ({row_reg, col_reg}<19'b0110001100011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0110001100011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0110001100011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0110001100011101010) && ({row_reg, col_reg}<19'b0110001100011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110001100011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0110001100011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110001100011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0110001100011101111) && ({row_reg, col_reg}<19'b0110001100100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110001100100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0110001100100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0110001100100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0110001100100000100) && ({row_reg, col_reg}<19'b0110001100101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0110001100101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0110001100101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0110001100110000000) && ({row_reg, col_reg}<19'b0110001100110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110001100110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0110001100110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0110001100110011010) && ({row_reg, col_reg}<19'b0110001110011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0110001110011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0110001110011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0110001110011101010) && ({row_reg, col_reg}<19'b0110001110011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110001110011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0110001110011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110001110011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0110001110011101111) && ({row_reg, col_reg}<19'b0110001110100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110001110100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0110001110100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0110001110100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0110001110100000100) && ({row_reg, col_reg}<19'b0110001110101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0110001110101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0110001110101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0110001110110000000) && ({row_reg, col_reg}<19'b0110001110110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110001110110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0110001110110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0110001110110011010) && ({row_reg, col_reg}<19'b0110010000011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0110010000011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0110010000011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0110010000011101010) && ({row_reg, col_reg}<19'b0110010000011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110010000011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0110010000011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110010000011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0110010000011101111) && ({row_reg, col_reg}<19'b0110010000100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110010000100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0110010000100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0110010000100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0110010000100000100) && ({row_reg, col_reg}<19'b0110010000101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0110010000101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0110010000101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0110010000110000000) && ({row_reg, col_reg}<19'b0110010000110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110010000110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0110010000110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0110010000110011010) && ({row_reg, col_reg}<19'b0110010010011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0110010010011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0110010010011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0110010010011101010) && ({row_reg, col_reg}<19'b0110010010011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110010010011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0110010010011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110010010011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0110010010011101111) && ({row_reg, col_reg}<19'b0110010010100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110010010100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0110010010100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0110010010100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0110010010100000100) && ({row_reg, col_reg}<19'b0110010010101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0110010010101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0110010010101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0110010010110000000) && ({row_reg, col_reg}<19'b0110010010110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110010010110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0110010010110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0110010010110011010) && ({row_reg, col_reg}<19'b0110010100011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0110010100011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0110010100011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0110010100011101010) && ({row_reg, col_reg}<19'b0110010100011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110010100011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0110010100011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110010100011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0110010100011101111) && ({row_reg, col_reg}<19'b0110010100100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110010100100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0110010100100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0110010100100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0110010100100000100) && ({row_reg, col_reg}<19'b0110010100101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0110010100101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0110010100101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0110010100110000000) && ({row_reg, col_reg}<19'b0110010100110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110010100110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0110010100110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0110010100110011010) && ({row_reg, col_reg}<19'b0110010110011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0110010110011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0110010110011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0110010110011101010) && ({row_reg, col_reg}<19'b0110010110011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110010110011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0110010110011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110010110011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0110010110011101111) && ({row_reg, col_reg}<19'b0110010110100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110010110100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0110010110100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0110010110100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0110010110100000100) && ({row_reg, col_reg}<19'b0110010110101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0110010110101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0110010110101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0110010110110000000) && ({row_reg, col_reg}<19'b0110010110110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110010110110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0110010110110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0110010110110011010) && ({row_reg, col_reg}<19'b0110011000011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0110011000011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0110011000011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0110011000011101010) && ({row_reg, col_reg}<19'b0110011000011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110011000011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0110011000011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110011000011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0110011000011101111) && ({row_reg, col_reg}<19'b0110011000100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110011000100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0110011000100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0110011000100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0110011000100000100) && ({row_reg, col_reg}<19'b0110011000101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0110011000101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0110011000101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0110011000110000000) && ({row_reg, col_reg}<19'b0110011000110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110011000110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0110011000110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0110011000110011010) && ({row_reg, col_reg}<19'b0110011010011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0110011010011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0110011010011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0110011010011101010) && ({row_reg, col_reg}<19'b0110011010011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110011010011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0110011010011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110011010011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0110011010011101111) && ({row_reg, col_reg}<19'b0110011010100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110011010100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0110011010100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0110011010100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0110011010100000100) && ({row_reg, col_reg}<19'b0110011010101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0110011010101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0110011010101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0110011010110000000) && ({row_reg, col_reg}<19'b0110011010110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110011010110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0110011010110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0110011010110011010) && ({row_reg, col_reg}<19'b0110011100011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0110011100011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0110011100011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0110011100011101010) && ({row_reg, col_reg}<19'b0110011100011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110011100011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0110011100011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110011100011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0110011100011101111) && ({row_reg, col_reg}<19'b0110011100100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110011100100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0110011100100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0110011100100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0110011100100000100) && ({row_reg, col_reg}<19'b0110011100101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0110011100101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0110011100101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0110011100110000000) && ({row_reg, col_reg}<19'b0110011100110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110011100110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0110011100110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0110011100110011010) && ({row_reg, col_reg}<19'b0110011110011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0110011110011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0110011110011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0110011110011101010) && ({row_reg, col_reg}<19'b0110011110011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110011110011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0110011110011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110011110011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0110011110011101111) && ({row_reg, col_reg}<19'b0110011110100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110011110100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0110011110100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0110011110100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0110011110100000100) && ({row_reg, col_reg}<19'b0110011110101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0110011110101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0110011110101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0110011110110000000) && ({row_reg, col_reg}<19'b0110011110110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110011110110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0110011110110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0110011110110011010) && ({row_reg, col_reg}<19'b0110100000011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0110100000011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0110100000011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0110100000011101010) && ({row_reg, col_reg}<19'b0110100000011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110100000011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0110100000011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110100000011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0110100000011101111) && ({row_reg, col_reg}<19'b0110100000100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110100000100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0110100000100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0110100000100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0110100000100000100) && ({row_reg, col_reg}<19'b0110100000101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0110100000101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0110100000101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0110100000110000000) && ({row_reg, col_reg}<19'b0110100000110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110100000110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0110100000110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0110100000110011010) && ({row_reg, col_reg}<19'b0110100010011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0110100010011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0110100010011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0110100010011101010) && ({row_reg, col_reg}<19'b0110100010011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110100010011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0110100010011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110100010011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0110100010011101111) && ({row_reg, col_reg}<19'b0110100010100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110100010100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0110100010100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0110100010100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0110100010100000100) && ({row_reg, col_reg}<19'b0110100010101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0110100010101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0110100010101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0110100010110000000) && ({row_reg, col_reg}<19'b0110100010110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110100010110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0110100010110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0110100010110011010) && ({row_reg, col_reg}<19'b0110100100011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0110100100011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0110100100011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0110100100011101010) && ({row_reg, col_reg}<19'b0110100100011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110100100011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0110100100011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110100100011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0110100100011101111) && ({row_reg, col_reg}<19'b0110100100100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110100100100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0110100100100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0110100100100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0110100100100000100) && ({row_reg, col_reg}<19'b0110100100101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0110100100101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0110100100101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0110100100110000000) && ({row_reg, col_reg}<19'b0110100100110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110100100110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0110100100110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0110100100110011010) && ({row_reg, col_reg}<19'b0110100110011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0110100110011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0110100110011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0110100110011101010) && ({row_reg, col_reg}<19'b0110100110011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110100110011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0110100110011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110100110011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0110100110011101111) && ({row_reg, col_reg}<19'b0110100110100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110100110100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0110100110100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0110100110100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0110100110100000100) && ({row_reg, col_reg}<19'b0110100110101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0110100110101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0110100110101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0110100110110000000) && ({row_reg, col_reg}<19'b0110100110110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110100110110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0110100110110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0110100110110011010) && ({row_reg, col_reg}<19'b0110101000011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0110101000011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0110101000011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0110101000011101010) && ({row_reg, col_reg}<19'b0110101000011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110101000011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0110101000011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110101000011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0110101000011101111) && ({row_reg, col_reg}<19'b0110101000100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110101000100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0110101000100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0110101000100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0110101000100000100) && ({row_reg, col_reg}<19'b0110101000101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0110101000101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0110101000101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0110101000110000000) && ({row_reg, col_reg}<19'b0110101000110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110101000110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0110101000110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0110101000110011010) && ({row_reg, col_reg}<19'b0110101010011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0110101010011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0110101010011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0110101010011101010) && ({row_reg, col_reg}<19'b0110101010011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110101010011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0110101010011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110101010011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0110101010011101111) && ({row_reg, col_reg}<19'b0110101010100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110101010100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0110101010100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0110101010100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0110101010100000100) && ({row_reg, col_reg}<19'b0110101010101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0110101010101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0110101010101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0110101010110000000) && ({row_reg, col_reg}<19'b0110101010110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110101010110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0110101010110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0110101010110011010) && ({row_reg, col_reg}<19'b0110101100011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0110101100011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0110101100011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0110101100011101010) && ({row_reg, col_reg}<19'b0110101100011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110101100011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0110101100011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110101100011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0110101100011101111) && ({row_reg, col_reg}<19'b0110101100100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110101100100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0110101100100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0110101100100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0110101100100000100) && ({row_reg, col_reg}<19'b0110101100101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0110101100101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0110101100101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0110101100110000000) && ({row_reg, col_reg}<19'b0110101100110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110101100110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0110101100110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0110101100110011010) && ({row_reg, col_reg}<19'b0110101110011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0110101110011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0110101110011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0110101110011101010) && ({row_reg, col_reg}<19'b0110101110011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110101110011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0110101110011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110101110011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0110101110011101111) && ({row_reg, col_reg}<19'b0110101110100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110101110100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0110101110100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0110101110100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0110101110100000100) && ({row_reg, col_reg}<19'b0110101110101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0110101110101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0110101110101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0110101110110000000) && ({row_reg, col_reg}<19'b0110101110110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110101110110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0110101110110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0110101110110011010) && ({row_reg, col_reg}<19'b0110110000011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0110110000011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0110110000011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0110110000011101010) && ({row_reg, col_reg}<19'b0110110000011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110110000011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0110110000011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110110000011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0110110000011101111) && ({row_reg, col_reg}<19'b0110110000100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110110000100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0110110000100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0110110000100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0110110000100000100) && ({row_reg, col_reg}<19'b0110110000101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0110110000101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0110110000101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0110110000110000000) && ({row_reg, col_reg}<19'b0110110000110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110110000110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0110110000110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0110110000110011010) && ({row_reg, col_reg}<19'b0110110010011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0110110010011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0110110010011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0110110010011101010) && ({row_reg, col_reg}<19'b0110110010011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110110010011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0110110010011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110110010011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0110110010011101111) && ({row_reg, col_reg}<19'b0110110010100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110110010100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0110110010100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0110110010100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0110110010100000100) && ({row_reg, col_reg}<19'b0110110010101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0110110010101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0110110010101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0110110010110000000) && ({row_reg, col_reg}<19'b0110110010110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110110010110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0110110010110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0110110010110011010) && ({row_reg, col_reg}<19'b0110110100011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0110110100011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0110110100011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0110110100011101010) && ({row_reg, col_reg}<19'b0110110100011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110110100011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0110110100011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110110100011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0110110100011101111) && ({row_reg, col_reg}<19'b0110110100100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110110100100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0110110100100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0110110100100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0110110100100000100) && ({row_reg, col_reg}<19'b0110110100101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0110110100101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0110110100101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0110110100110000000) && ({row_reg, col_reg}<19'b0110110100110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110110100110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0110110100110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0110110100110011010) && ({row_reg, col_reg}<19'b0110110110011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0110110110011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0110110110011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0110110110011101010) && ({row_reg, col_reg}<19'b0110110110011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110110110011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0110110110011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110110110011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0110110110011101111) && ({row_reg, col_reg}<19'b0110110110100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110110110100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0110110110100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0110110110100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0110110110100000100) && ({row_reg, col_reg}<19'b0110110110101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0110110110101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0110110110101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0110110110110000000) && ({row_reg, col_reg}<19'b0110110110110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110110110110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0110110110110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0110110110110011010) && ({row_reg, col_reg}<19'b0110111000011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0110111000011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0110111000011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0110111000011101010) && ({row_reg, col_reg}<19'b0110111000011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110111000011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0110111000011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110111000011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0110111000011101111) && ({row_reg, col_reg}<19'b0110111000100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110111000100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0110111000100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0110111000100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0110111000100000100) && ({row_reg, col_reg}<19'b0110111000101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0110111000101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0110111000101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0110111000110000000) && ({row_reg, col_reg}<19'b0110111000110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110111000110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0110111000110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0110111000110011010) && ({row_reg, col_reg}<19'b0110111010011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0110111010011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0110111010011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0110111010011101010) && ({row_reg, col_reg}<19'b0110111010011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110111010011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0110111010011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110111010011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0110111010011101111) && ({row_reg, col_reg}<19'b0110111010100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110111010100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0110111010100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0110111010100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0110111010100000100) && ({row_reg, col_reg}<19'b0110111010101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0110111010101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0110111010101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0110111010110000000) && ({row_reg, col_reg}<19'b0110111010110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110111010110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0110111010110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0110111010110011010) && ({row_reg, col_reg}<19'b0110111100011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0110111100011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0110111100011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0110111100011101010) && ({row_reg, col_reg}<19'b0110111100011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110111100011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0110111100011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110111100011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0110111100011101111) && ({row_reg, col_reg}<19'b0110111100100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110111100100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0110111100100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0110111100100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0110111100100000100) && ({row_reg, col_reg}<19'b0110111100101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0110111100101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0110111100101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0110111100110000000) && ({row_reg, col_reg}<19'b0110111100110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110111100110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0110111100110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0110111100110011010) && ({row_reg, col_reg}<19'b0110111110011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0110111110011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0110111110011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0110111110011101010) && ({row_reg, col_reg}<19'b0110111110011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110111110011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0110111110011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110111110011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0110111110011101111) && ({row_reg, col_reg}<19'b0110111110100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110111110100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0110111110100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0110111110100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0110111110100000100) && ({row_reg, col_reg}<19'b0110111110101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0110111110101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0110111110101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0110111110110000000) && ({row_reg, col_reg}<19'b0110111110110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110111110110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0110111110110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0110111110110011010) && ({row_reg, col_reg}<19'b0111000000011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111000000011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0111000000011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111000000011101010) && ({row_reg, col_reg}<19'b0111000000011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111000000011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0111000000011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111000000011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111000000011101111) && ({row_reg, col_reg}<19'b0111000000100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111000000100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0111000000100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0111000000100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0111000000100000100) && ({row_reg, col_reg}<19'b0111000000101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111000000101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0111000000101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111000000110000000) && ({row_reg, col_reg}<19'b0111000000110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111000000110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0111000000110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0111000000110011010) && ({row_reg, col_reg}<19'b0111000010011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111000010011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0111000010011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111000010011101010) && ({row_reg, col_reg}<19'b0111000010011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111000010011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0111000010011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111000010011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111000010011101111) && ({row_reg, col_reg}<19'b0111000010100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111000010100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0111000010100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0111000010100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0111000010100000100) && ({row_reg, col_reg}<19'b0111000010101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111000010101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0111000010101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111000010110000000) && ({row_reg, col_reg}<19'b0111000010110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111000010110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0111000010110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0111000010110011010) && ({row_reg, col_reg}<19'b0111000100011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111000100011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0111000100011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111000100011101010) && ({row_reg, col_reg}<19'b0111000100011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111000100011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0111000100011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111000100011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111000100011101111) && ({row_reg, col_reg}<19'b0111000100100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111000100100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0111000100100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0111000100100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0111000100100000100) && ({row_reg, col_reg}<19'b0111000100101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111000100101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0111000100101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111000100110000000) && ({row_reg, col_reg}<19'b0111000100110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111000100110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0111000100110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0111000100110011010) && ({row_reg, col_reg}<19'b0111000110011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111000110011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0111000110011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111000110011101010) && ({row_reg, col_reg}<19'b0111000110011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111000110011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0111000110011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111000110011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111000110011101111) && ({row_reg, col_reg}<19'b0111000110100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111000110100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0111000110100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0111000110100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0111000110100000100) && ({row_reg, col_reg}<19'b0111000110101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111000110101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0111000110101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111000110110000000) && ({row_reg, col_reg}<19'b0111000110110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111000110110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0111000110110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0111000110110011010) && ({row_reg, col_reg}<19'b0111001000011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111001000011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0111001000011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111001000011101010) && ({row_reg, col_reg}<19'b0111001000011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111001000011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0111001000011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111001000011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111001000011101111) && ({row_reg, col_reg}<19'b0111001000100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111001000100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0111001000100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0111001000100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0111001000100000100) && ({row_reg, col_reg}<19'b0111001000101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111001000101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0111001000101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111001000110000000) && ({row_reg, col_reg}<19'b0111001000110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111001000110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0111001000110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0111001000110011010) && ({row_reg, col_reg}<19'b0111001010011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111001010011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0111001010011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111001010011101010) && ({row_reg, col_reg}<19'b0111001010011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111001010011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0111001010011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111001010011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111001010011101111) && ({row_reg, col_reg}<19'b0111001010100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111001010100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0111001010100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0111001010100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0111001010100000100) && ({row_reg, col_reg}<19'b0111001010101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111001010101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0111001010101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111001010110000000) && ({row_reg, col_reg}<19'b0111001010110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111001010110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0111001010110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0111001010110011010) && ({row_reg, col_reg}<19'b0111001100011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111001100011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0111001100011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111001100011101010) && ({row_reg, col_reg}<19'b0111001100011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111001100011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0111001100011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111001100011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111001100011101111) && ({row_reg, col_reg}<19'b0111001100100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111001100100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0111001100100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0111001100100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0111001100100000100) && ({row_reg, col_reg}<19'b0111001100101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111001100101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0111001100101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111001100110000000) && ({row_reg, col_reg}<19'b0111001100110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111001100110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0111001100110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0111001100110011010) && ({row_reg, col_reg}<19'b0111001110011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111001110011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0111001110011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111001110011101010) && ({row_reg, col_reg}<19'b0111001110011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111001110011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0111001110011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111001110011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111001110011101111) && ({row_reg, col_reg}<19'b0111001110100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111001110100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0111001110100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0111001110100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0111001110100000100) && ({row_reg, col_reg}<19'b0111001110101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111001110101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0111001110101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111001110110000000) && ({row_reg, col_reg}<19'b0111001110110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111001110110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0111001110110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0111001110110011010) && ({row_reg, col_reg}<19'b0111010000011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111010000011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0111010000011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111010000011101010) && ({row_reg, col_reg}<19'b0111010000011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111010000011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0111010000011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111010000011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111010000011101111) && ({row_reg, col_reg}<19'b0111010000100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111010000100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0111010000100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0111010000100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0111010000100000100) && ({row_reg, col_reg}<19'b0111010000101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111010000101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0111010000101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111010000110000000) && ({row_reg, col_reg}<19'b0111010000110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111010000110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0111010000110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0111010000110011010) && ({row_reg, col_reg}<19'b0111010010011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111010010011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0111010010011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111010010011101010) && ({row_reg, col_reg}<19'b0111010010011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111010010011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0111010010011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111010010011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111010010011101111) && ({row_reg, col_reg}<19'b0111010010100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111010010100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0111010010100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0111010010100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0111010010100000100) && ({row_reg, col_reg}<19'b0111010010101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111010010101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0111010010101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111010010110000000) && ({row_reg, col_reg}<19'b0111010010110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111010010110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0111010010110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0111010010110011010) && ({row_reg, col_reg}<19'b0111010100011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111010100011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0111010100011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111010100011101010) && ({row_reg, col_reg}<19'b0111010100011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111010100011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0111010100011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111010100011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111010100011101111) && ({row_reg, col_reg}<19'b0111010100100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111010100100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0111010100100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0111010100100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0111010100100000100) && ({row_reg, col_reg}<19'b0111010100101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111010100101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0111010100101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111010100110000000) && ({row_reg, col_reg}<19'b0111010100110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111010100110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0111010100110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0111010100110011010) && ({row_reg, col_reg}<19'b0111010110011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111010110011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0111010110011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111010110011101010) && ({row_reg, col_reg}<19'b0111010110011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111010110011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0111010110011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111010110011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111010110011101111) && ({row_reg, col_reg}<19'b0111010110100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111010110100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0111010110100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0111010110100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0111010110100000100) && ({row_reg, col_reg}<19'b0111010110101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111010110101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0111010110101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111010110110000000) && ({row_reg, col_reg}<19'b0111010110110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111010110110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0111010110110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0111010110110011010) && ({row_reg, col_reg}<19'b0111011000011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111011000011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0111011000011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111011000011101010) && ({row_reg, col_reg}<19'b0111011000011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111011000011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0111011000011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111011000011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111011000011101111) && ({row_reg, col_reg}<19'b0111011000100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111011000100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0111011000100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0111011000100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0111011000100000100) && ({row_reg, col_reg}<19'b0111011000101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111011000101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0111011000101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111011000110000000) && ({row_reg, col_reg}<19'b0111011000110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111011000110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0111011000110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0111011000110011010) && ({row_reg, col_reg}<19'b0111011010011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111011010011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0111011010011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111011010011101010) && ({row_reg, col_reg}<19'b0111011010011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111011010011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0111011010011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111011010011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111011010011101111) && ({row_reg, col_reg}<19'b0111011010100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111011010100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0111011010100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0111011010100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0111011010100000100) && ({row_reg, col_reg}<19'b0111011010101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111011010101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0111011010101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111011010110000000) && ({row_reg, col_reg}<19'b0111011010110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111011010110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0111011010110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0111011010110011010) && ({row_reg, col_reg}<19'b0111011100011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111011100011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0111011100011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111011100011101010) && ({row_reg, col_reg}<19'b0111011100011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111011100011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0111011100011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111011100011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111011100011101111) && ({row_reg, col_reg}<19'b0111011100100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111011100100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0111011100100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0111011100100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0111011100100000100) && ({row_reg, col_reg}<19'b0111011100101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111011100101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0111011100101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111011100110000000) && ({row_reg, col_reg}<19'b0111011100110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111011100110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0111011100110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0111011100110011010) && ({row_reg, col_reg}<19'b0111011110011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111011110011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0111011110011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111011110011101010) && ({row_reg, col_reg}<19'b0111011110011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111011110011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0111011110011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111011110011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111011110011101111) && ({row_reg, col_reg}<19'b0111011110100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111011110100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0111011110100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0111011110100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0111011110100000100) && ({row_reg, col_reg}<19'b0111011110101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111011110101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0111011110101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111011110110000000) && ({row_reg, col_reg}<19'b0111011110110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111011110110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0111011110110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0111011110110011010) && ({row_reg, col_reg}<19'b0111100000011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111100000011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0111100000011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111100000011101010) && ({row_reg, col_reg}<19'b0111100000011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111100000011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0111100000011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111100000011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111100000011101111) && ({row_reg, col_reg}<19'b0111100000100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111100000100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0111100000100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0111100000100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0111100000100000100) && ({row_reg, col_reg}<19'b0111100000101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111100000101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0111100000101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111100000110000000) && ({row_reg, col_reg}<19'b0111100000110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111100000110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0111100000110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0111100000110011010) && ({row_reg, col_reg}<19'b0111100010011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111100010011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0111100010011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111100010011101010) && ({row_reg, col_reg}<19'b0111100010011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111100010011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0111100010011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111100010011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111100010011101111) && ({row_reg, col_reg}<19'b0111100010100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111100010100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0111100010100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0111100010100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0111100010100000100) && ({row_reg, col_reg}<19'b0111100010101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111100010101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0111100010101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111100010110000000) && ({row_reg, col_reg}<19'b0111100010110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111100010110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0111100010110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0111100010110011010) && ({row_reg, col_reg}<19'b0111100100011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111100100011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0111100100011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111100100011101010) && ({row_reg, col_reg}<19'b0111100100011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111100100011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0111100100011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111100100011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111100100011101111) && ({row_reg, col_reg}<19'b0111100100100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111100100100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0111100100100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0111100100100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0111100100100000100) && ({row_reg, col_reg}<19'b0111100100101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111100100101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0111100100101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111100100110000000) && ({row_reg, col_reg}<19'b0111100100110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111100100110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0111100100110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0111100100110011010) && ({row_reg, col_reg}<19'b0111100110011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111100110011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0111100110011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111100110011101010) && ({row_reg, col_reg}<19'b0111100110011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111100110011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0111100110011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111100110011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111100110011101111) && ({row_reg, col_reg}<19'b0111100110100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111100110100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0111100110100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0111100110100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0111100110100000100) && ({row_reg, col_reg}<19'b0111100110101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111100110101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0111100110101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111100110110000000) && ({row_reg, col_reg}<19'b0111100110110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111100110110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0111100110110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0111100110110011010) && ({row_reg, col_reg}<19'b0111101000011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111101000011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0111101000011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111101000011101010) && ({row_reg, col_reg}<19'b0111101000011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111101000011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0111101000011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111101000011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111101000011101111) && ({row_reg, col_reg}<19'b0111101000100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111101000100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0111101000100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0111101000100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0111101000100000100) && ({row_reg, col_reg}<19'b0111101000101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111101000101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0111101000101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111101000110000000) && ({row_reg, col_reg}<19'b0111101000110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111101000110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0111101000110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0111101000110011010) && ({row_reg, col_reg}<19'b0111101010011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111101010011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0111101010011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111101010011101010) && ({row_reg, col_reg}<19'b0111101010011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111101010011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0111101010011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111101010011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111101010011101111) && ({row_reg, col_reg}<19'b0111101010100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111101010100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0111101010100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0111101010100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0111101010100000100) && ({row_reg, col_reg}<19'b0111101010101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111101010101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0111101010101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111101010110000000) && ({row_reg, col_reg}<19'b0111101010110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111101010110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0111101010110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0111101010110011010) && ({row_reg, col_reg}<19'b0111101100011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111101100011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0111101100011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111101100011101010) && ({row_reg, col_reg}<19'b0111101100011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111101100011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0111101100011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111101100011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111101100011101111) && ({row_reg, col_reg}<19'b0111101100100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111101100100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0111101100100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0111101100100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0111101100100000100) && ({row_reg, col_reg}<19'b0111101100101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111101100101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0111101100101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111101100110000000) && ({row_reg, col_reg}<19'b0111101100110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111101100110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0111101100110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0111101100110011010) && ({row_reg, col_reg}<19'b0111101110011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111101110011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0111101110011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111101110011101010) && ({row_reg, col_reg}<19'b0111101110011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111101110011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0111101110011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111101110011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111101110011101111) && ({row_reg, col_reg}<19'b0111101110100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111101110100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0111101110100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0111101110100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0111101110100000100) && ({row_reg, col_reg}<19'b0111101110101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111101110101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0111101110101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111101110110000000) && ({row_reg, col_reg}<19'b0111101110110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111101110110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0111101110110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0111101110110011010) && ({row_reg, col_reg}<19'b0111110000011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111110000011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0111110000011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111110000011101010) && ({row_reg, col_reg}<19'b0111110000011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111110000011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0111110000011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111110000011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111110000011101111) && ({row_reg, col_reg}<19'b0111110000100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111110000100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0111110000100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0111110000100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0111110000100000100) && ({row_reg, col_reg}<19'b0111110000101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111110000101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0111110000101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111110000110000000) && ({row_reg, col_reg}<19'b0111110000110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111110000110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0111110000110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0111110000110011010) && ({row_reg, col_reg}<19'b0111110010011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111110010011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0111110010011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111110010011101010) && ({row_reg, col_reg}<19'b0111110010011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111110010011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0111110010011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111110010011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111110010011101111) && ({row_reg, col_reg}<19'b0111110010100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111110010100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0111110010100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0111110010100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0111110010100000100) && ({row_reg, col_reg}<19'b0111110010101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111110010101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0111110010101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111110010110000000) && ({row_reg, col_reg}<19'b0111110010110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111110010110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0111110010110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0111110010110011010) && ({row_reg, col_reg}<19'b0111110100011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111110100011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0111110100011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111110100011101010) && ({row_reg, col_reg}<19'b0111110100011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111110100011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0111110100011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111110100011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111110100011101111) && ({row_reg, col_reg}<19'b0111110100100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111110100100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0111110100100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0111110100100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0111110100100000100) && ({row_reg, col_reg}<19'b0111110100101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111110100101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0111110100101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111110100110000000) && ({row_reg, col_reg}<19'b0111110100110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111110100110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0111110100110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0111110100110011010) && ({row_reg, col_reg}<19'b0111110110011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111110110011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0111110110011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111110110011101010) && ({row_reg, col_reg}<19'b0111110110011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111110110011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0111110110011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111110110011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111110110011101111) && ({row_reg, col_reg}<19'b0111110110100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111110110100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0111110110100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0111110110100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0111110110100000100) && ({row_reg, col_reg}<19'b0111110110101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111110110101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0111110110101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111110110110000000) && ({row_reg, col_reg}<19'b0111110110110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111110110110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0111110110110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0111110110110011010) && ({row_reg, col_reg}<19'b0111111000011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111111000011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0111111000011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111111000011101010) && ({row_reg, col_reg}<19'b0111111000011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111111000011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0111111000011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111111000011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111111000011101111) && ({row_reg, col_reg}<19'b0111111000100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111111000100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0111111000100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0111111000100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0111111000100000100) && ({row_reg, col_reg}<19'b0111111000101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111111000101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0111111000101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111111000110000000) && ({row_reg, col_reg}<19'b0111111000110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111111000110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0111111000110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0111111000110011010) && ({row_reg, col_reg}<19'b0111111010011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111111010011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0111111010011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111111010011101010) && ({row_reg, col_reg}<19'b0111111010011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111111010011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0111111010011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111111010011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111111010011101111) && ({row_reg, col_reg}<19'b0111111010100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111111010100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0111111010100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0111111010100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0111111010100000100) && ({row_reg, col_reg}<19'b0111111010101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111111010101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0111111010101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111111010110000000) && ({row_reg, col_reg}<19'b0111111010110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111111010110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0111111010110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0111111010110011010) && ({row_reg, col_reg}<19'b0111111100011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111111100011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0111111100011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111111100011101010) && ({row_reg, col_reg}<19'b0111111100011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111111100011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0111111100011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111111100011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111111100011101111) && ({row_reg, col_reg}<19'b0111111100100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111111100100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0111111100100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0111111100100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0111111100100000100) && ({row_reg, col_reg}<19'b0111111100101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111111100101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0111111100101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111111100110000000) && ({row_reg, col_reg}<19'b0111111100110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111111100110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0111111100110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0111111100110011010) && ({row_reg, col_reg}<19'b0111111110011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111111110011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0111111110011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111111110011101010) && ({row_reg, col_reg}<19'b0111111110011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111111110011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0111111110011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111111110011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111111110011101111) && ({row_reg, col_reg}<19'b0111111110100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111111110100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0111111110100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0111111110100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0111111110100000100) && ({row_reg, col_reg}<19'b0111111110101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111111110101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0111111110101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111111110110000000) && ({row_reg, col_reg}<19'b0111111110110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111111110110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0111111110110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0111111110110011010) && ({row_reg, col_reg}<19'b1000000000011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000000000011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1000000000011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000000000011101010) && ({row_reg, col_reg}<19'b1000000000011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000000000011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1000000000011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000000000011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000000000011101111) && ({row_reg, col_reg}<19'b1000000000100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000000000100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1000000000100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1000000000100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1000000000100000100) && ({row_reg, col_reg}<19'b1000000000101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000000000101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1000000000101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000000000110000000) && ({row_reg, col_reg}<19'b1000000000110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000000000110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1000000000110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1000000000110011010) && ({row_reg, col_reg}<19'b1000000010011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000000010011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1000000010011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000000010011101010) && ({row_reg, col_reg}<19'b1000000010011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000000010011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1000000010011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000000010011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000000010011101111) && ({row_reg, col_reg}<19'b1000000010100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000000010100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1000000010100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1000000010100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1000000010100000100) && ({row_reg, col_reg}<19'b1000000010101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000000010101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1000000010101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000000010110000000) && ({row_reg, col_reg}<19'b1000000010110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000000010110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1000000010110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1000000010110011010) && ({row_reg, col_reg}<19'b1000000100011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000000100011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1000000100011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000000100011101010) && ({row_reg, col_reg}<19'b1000000100011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000000100011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1000000100011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000000100011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000000100011101111) && ({row_reg, col_reg}<19'b1000000100100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000000100100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1000000100100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1000000100100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1000000100100000100) && ({row_reg, col_reg}<19'b1000000100101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000000100101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1000000100101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000000100110000000) && ({row_reg, col_reg}<19'b1000000100110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000000100110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1000000100110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1000000100110011010) && ({row_reg, col_reg}<19'b1000000110011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000000110011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1000000110011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000000110011101010) && ({row_reg, col_reg}<19'b1000000110011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000000110011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1000000110011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000000110011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000000110011101111) && ({row_reg, col_reg}<19'b1000000110100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000000110100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1000000110100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1000000110100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1000000110100000100) && ({row_reg, col_reg}<19'b1000000110101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000000110101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1000000110101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000000110110000000) && ({row_reg, col_reg}<19'b1000000110110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000000110110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1000000110110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1000000110110011010) && ({row_reg, col_reg}<19'b1000001000011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000001000011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1000001000011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000001000011101010) && ({row_reg, col_reg}<19'b1000001000011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000001000011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1000001000011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000001000011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000001000011101111) && ({row_reg, col_reg}<19'b1000001000100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000001000100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1000001000100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1000001000100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1000001000100000100) && ({row_reg, col_reg}<19'b1000001000101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000001000101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1000001000101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000001000110000000) && ({row_reg, col_reg}<19'b1000001000110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000001000110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1000001000110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1000001000110011010) && ({row_reg, col_reg}<19'b1000001010011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000001010011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1000001010011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000001010011101010) && ({row_reg, col_reg}<19'b1000001010011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000001010011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1000001010011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000001010011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000001010011101111) && ({row_reg, col_reg}<19'b1000001010100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000001010100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1000001010100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1000001010100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1000001010100000100) && ({row_reg, col_reg}<19'b1000001010101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000001010101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1000001010101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000001010110000000) && ({row_reg, col_reg}<19'b1000001010110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000001010110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1000001010110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1000001010110011010) && ({row_reg, col_reg}<19'b1000001100011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000001100011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1000001100011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000001100011101010) && ({row_reg, col_reg}<19'b1000001100011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000001100011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1000001100011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000001100011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000001100011101111) && ({row_reg, col_reg}<19'b1000001100100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000001100100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1000001100100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1000001100100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1000001100100000100) && ({row_reg, col_reg}<19'b1000001100101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000001100101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1000001100101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000001100110000000) && ({row_reg, col_reg}<19'b1000001100110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000001100110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1000001100110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1000001100110011010) && ({row_reg, col_reg}<19'b1000001110011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000001110011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1000001110011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000001110011101010) && ({row_reg, col_reg}<19'b1000001110011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000001110011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1000001110011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000001110011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000001110011101111) && ({row_reg, col_reg}<19'b1000001110100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000001110100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1000001110100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1000001110100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1000001110100000100) && ({row_reg, col_reg}<19'b1000001110101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000001110101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1000001110101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000001110110000000) && ({row_reg, col_reg}<19'b1000001110110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000001110110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1000001110110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1000001110110011010) && ({row_reg, col_reg}<19'b1000010000011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000010000011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1000010000011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000010000011101010) && ({row_reg, col_reg}<19'b1000010000011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000010000011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1000010000011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000010000011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000010000011101111) && ({row_reg, col_reg}<19'b1000010000100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000010000100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1000010000100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1000010000100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1000010000100000100) && ({row_reg, col_reg}<19'b1000010000101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000010000101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1000010000101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000010000110000000) && ({row_reg, col_reg}<19'b1000010000110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000010000110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1000010000110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1000010000110011010) && ({row_reg, col_reg}<19'b1000010010011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000010010011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1000010010011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000010010011101010) && ({row_reg, col_reg}<19'b1000010010011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000010010011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1000010010011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000010010011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000010010011101111) && ({row_reg, col_reg}<19'b1000010010100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000010010100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1000010010100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1000010010100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1000010010100000100) && ({row_reg, col_reg}<19'b1000010010101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000010010101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1000010010101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000010010110000000) && ({row_reg, col_reg}<19'b1000010010110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000010010110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1000010010110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1000010010110011010) && ({row_reg, col_reg}<19'b1000010100011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000010100011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1000010100011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000010100011101010) && ({row_reg, col_reg}<19'b1000010100011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000010100011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1000010100011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000010100011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000010100011101111) && ({row_reg, col_reg}<19'b1000010100100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000010100100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1000010100100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1000010100100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1000010100100000100) && ({row_reg, col_reg}<19'b1000010100101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000010100101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1000010100101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000010100110000000) && ({row_reg, col_reg}<19'b1000010100110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000010100110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1000010100110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1000010100110011010) && ({row_reg, col_reg}<19'b1000010110011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000010110011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1000010110011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000010110011101010) && ({row_reg, col_reg}<19'b1000010110011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000010110011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1000010110011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000010110011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000010110011101111) && ({row_reg, col_reg}<19'b1000010110100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000010110100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1000010110100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1000010110100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1000010110100000100) && ({row_reg, col_reg}<19'b1000010110101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000010110101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1000010110101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000010110110000000) && ({row_reg, col_reg}<19'b1000010110110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000010110110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1000010110110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1000010110110011010) && ({row_reg, col_reg}<19'b1000011000011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000011000011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1000011000011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000011000011101010) && ({row_reg, col_reg}<19'b1000011000011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000011000011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1000011000011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000011000011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000011000011101111) && ({row_reg, col_reg}<19'b1000011000100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000011000100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1000011000100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1000011000100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1000011000100000100) && ({row_reg, col_reg}<19'b1000011000101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000011000101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1000011000101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000011000110000000) && ({row_reg, col_reg}<19'b1000011000110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000011000110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1000011000110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1000011000110011010) && ({row_reg, col_reg}<19'b1000011010011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000011010011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1000011010011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000011010011101010) && ({row_reg, col_reg}<19'b1000011010011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000011010011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1000011010011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000011010011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000011010011101111) && ({row_reg, col_reg}<19'b1000011010100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000011010100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1000011010100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1000011010100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1000011010100000100) && ({row_reg, col_reg}<19'b1000011010101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000011010101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1000011010101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000011010110000000) && ({row_reg, col_reg}<19'b1000011010110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000011010110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1000011010110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1000011010110011010) && ({row_reg, col_reg}<19'b1000011100011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000011100011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1000011100011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000011100011101010) && ({row_reg, col_reg}<19'b1000011100011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000011100011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1000011100011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000011100011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000011100011101111) && ({row_reg, col_reg}<19'b1000011100100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000011100100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1000011100100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1000011100100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1000011100100000100) && ({row_reg, col_reg}<19'b1000011100101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000011100101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1000011100101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000011100110000000) && ({row_reg, col_reg}<19'b1000011100110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000011100110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1000011100110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1000011100110011010) && ({row_reg, col_reg}<19'b1000011110011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000011110011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1000011110011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000011110011101010) && ({row_reg, col_reg}<19'b1000011110011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000011110011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1000011110011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000011110011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000011110011101111) && ({row_reg, col_reg}<19'b1000011110100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000011110100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1000011110100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1000011110100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1000011110100000100) && ({row_reg, col_reg}<19'b1000011110101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000011110101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1000011110101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000011110110000000) && ({row_reg, col_reg}<19'b1000011110110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000011110110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1000011110110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1000011110110011010) && ({row_reg, col_reg}<19'b1000100000011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000100000011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1000100000011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000100000011101010) && ({row_reg, col_reg}<19'b1000100000011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000100000011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1000100000011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000100000011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000100000011101111) && ({row_reg, col_reg}<19'b1000100000100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000100000100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1000100000100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1000100000100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1000100000100000100) && ({row_reg, col_reg}<19'b1000100000101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000100000101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1000100000101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000100000110000000) && ({row_reg, col_reg}<19'b1000100000110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000100000110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1000100000110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1000100000110011010) && ({row_reg, col_reg}<19'b1000100010011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000100010011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1000100010011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000100010011101010) && ({row_reg, col_reg}<19'b1000100010011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000100010011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1000100010011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000100010011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000100010011101111) && ({row_reg, col_reg}<19'b1000100010100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000100010100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1000100010100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1000100010100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1000100010100000100) && ({row_reg, col_reg}<19'b1000100010101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000100010101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1000100010101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000100010110000000) && ({row_reg, col_reg}<19'b1000100010110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000100010110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1000100010110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1000100010110011010) && ({row_reg, col_reg}<19'b1000100100011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000100100011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1000100100011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000100100011101010) && ({row_reg, col_reg}<19'b1000100100011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000100100011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1000100100011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000100100011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000100100011101111) && ({row_reg, col_reg}<19'b1000100100100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000100100100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1000100100100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1000100100100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1000100100100000100) && ({row_reg, col_reg}<19'b1000100100101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000100100101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1000100100101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000100100110000000) && ({row_reg, col_reg}<19'b1000100100110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000100100110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1000100100110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1000100100110011010) && ({row_reg, col_reg}<19'b1000100110011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000100110011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1000100110011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000100110011101010) && ({row_reg, col_reg}<19'b1000100110011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000100110011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1000100110011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000100110011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000100110011101111) && ({row_reg, col_reg}<19'b1000100110100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000100110100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1000100110100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1000100110100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1000100110100000100) && ({row_reg, col_reg}<19'b1000100110101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000100110101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1000100110101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000100110110000000) && ({row_reg, col_reg}<19'b1000100110110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000100110110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1000100110110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1000100110110011010) && ({row_reg, col_reg}<19'b1000101000011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000101000011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1000101000011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000101000011101010) && ({row_reg, col_reg}<19'b1000101000011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000101000011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1000101000011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000101000011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000101000011101111) && ({row_reg, col_reg}<19'b1000101000100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000101000100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1000101000100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1000101000100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1000101000100000100) && ({row_reg, col_reg}<19'b1000101000101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000101000101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1000101000101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000101000110000000) && ({row_reg, col_reg}<19'b1000101000110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000101000110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1000101000110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1000101000110011010) && ({row_reg, col_reg}<19'b1000101010011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000101010011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1000101010011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000101010011101010) && ({row_reg, col_reg}<19'b1000101010011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000101010011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1000101010011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000101010011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000101010011101111) && ({row_reg, col_reg}<19'b1000101010100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000101010100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1000101010100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1000101010100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1000101010100000100) && ({row_reg, col_reg}<19'b1000101010101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000101010101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1000101010101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000101010110000000) && ({row_reg, col_reg}<19'b1000101010110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000101010110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1000101010110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1000101010110011010) && ({row_reg, col_reg}<19'b1000101100011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000101100011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1000101100011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000101100011101010) && ({row_reg, col_reg}<19'b1000101100011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000101100011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1000101100011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000101100011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000101100011101111) && ({row_reg, col_reg}<19'b1000101100100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000101100100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1000101100100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1000101100100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1000101100100000100) && ({row_reg, col_reg}<19'b1000101100101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000101100101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1000101100101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000101100110000000) && ({row_reg, col_reg}<19'b1000101100110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000101100110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1000101100110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1000101100110011010) && ({row_reg, col_reg}<19'b1000101110011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000101110011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1000101110011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000101110011101010) && ({row_reg, col_reg}<19'b1000101110011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000101110011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1000101110011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000101110011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000101110011101111) && ({row_reg, col_reg}<19'b1000101110100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000101110100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1000101110100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1000101110100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1000101110100000100) && ({row_reg, col_reg}<19'b1000101110101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000101110101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1000101110101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000101110110000000) && ({row_reg, col_reg}<19'b1000101110110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000101110110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1000101110110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1000101110110011010) && ({row_reg, col_reg}<19'b1000110000011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000110000011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1000110000011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000110000011101010) && ({row_reg, col_reg}<19'b1000110000011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000110000011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1000110000011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000110000011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000110000011101111) && ({row_reg, col_reg}<19'b1000110000100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000110000100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1000110000100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1000110000100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1000110000100000100) && ({row_reg, col_reg}<19'b1000110000101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000110000101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1000110000101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000110000110000000) && ({row_reg, col_reg}<19'b1000110000110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000110000110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1000110000110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1000110000110011010) && ({row_reg, col_reg}<19'b1000110010011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000110010011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1000110010011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000110010011101010) && ({row_reg, col_reg}<19'b1000110010011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000110010011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1000110010011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000110010011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000110010011101111) && ({row_reg, col_reg}<19'b1000110010100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000110010100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1000110010100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1000110010100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1000110010100000100) && ({row_reg, col_reg}<19'b1000110010101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000110010101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1000110010101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000110010110000000) && ({row_reg, col_reg}<19'b1000110010110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000110010110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1000110010110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1000110010110011010) && ({row_reg, col_reg}<19'b1000110100011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000110100011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1000110100011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000110100011101010) && ({row_reg, col_reg}<19'b1000110100011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000110100011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1000110100011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000110100011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000110100011101111) && ({row_reg, col_reg}<19'b1000110100100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000110100100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1000110100100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1000110100100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1000110100100000100) && ({row_reg, col_reg}<19'b1000110100101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000110100101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1000110100101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000110100110000000) && ({row_reg, col_reg}<19'b1000110100110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000110100110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1000110100110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1000110100110011010) && ({row_reg, col_reg}<19'b1000110110011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000110110011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1000110110011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000110110011101010) && ({row_reg, col_reg}<19'b1000110110011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000110110011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1000110110011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000110110011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000110110011101111) && ({row_reg, col_reg}<19'b1000110110100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000110110100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1000110110100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1000110110100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1000110110100000100) && ({row_reg, col_reg}<19'b1000110110101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000110110101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1000110110101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000110110110000000) && ({row_reg, col_reg}<19'b1000110110110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000110110110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1000110110110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1000110110110011010) && ({row_reg, col_reg}<19'b1000111000011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000111000011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1000111000011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000111000011101010) && ({row_reg, col_reg}<19'b1000111000011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000111000011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1000111000011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000111000011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000111000011101111) && ({row_reg, col_reg}<19'b1000111000100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000111000100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1000111000100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1000111000100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1000111000100000100) && ({row_reg, col_reg}<19'b1000111000101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000111000101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1000111000101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000111000110000000) && ({row_reg, col_reg}<19'b1000111000110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000111000110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1000111000110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1000111000110011010) && ({row_reg, col_reg}<19'b1000111010011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000111010011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1000111010011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000111010011101010) && ({row_reg, col_reg}<19'b1000111010011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000111010011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1000111010011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000111010011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000111010011101111) && ({row_reg, col_reg}<19'b1000111010100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000111010100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1000111010100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1000111010100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1000111010100000100) && ({row_reg, col_reg}<19'b1000111010101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000111010101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1000111010101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000111010110000000) && ({row_reg, col_reg}<19'b1000111010110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000111010110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1000111010110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1000111010110011010) && ({row_reg, col_reg}<19'b1000111100011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000111100011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1000111100011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000111100011101010) && ({row_reg, col_reg}<19'b1000111100011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000111100011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1000111100011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000111100011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000111100011101111) && ({row_reg, col_reg}<19'b1000111100100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000111100100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1000111100100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1000111100100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1000111100100000100) && ({row_reg, col_reg}<19'b1000111100101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000111100101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1000111100101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000111100110000000) && ({row_reg, col_reg}<19'b1000111100110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000111100110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1000111100110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1000111100110011010) && ({row_reg, col_reg}<19'b1000111110011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000111110011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1000111110011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000111110011101010) && ({row_reg, col_reg}<19'b1000111110011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000111110011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1000111110011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000111110011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000111110011101111) && ({row_reg, col_reg}<19'b1000111110100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000111110100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1000111110100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1000111110100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1000111110100000100) && ({row_reg, col_reg}<19'b1000111110101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000111110101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1000111110101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000111110110000000) && ({row_reg, col_reg}<19'b1000111110110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000111110110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1000111110110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1000111110110011010) && ({row_reg, col_reg}<19'b1001000000011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1001000000011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1001000000011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001000000011101010) && ({row_reg, col_reg}<19'b1001000000011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001000000011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1001000000011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001000000011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001000000011101111) && ({row_reg, col_reg}<19'b1001000000100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001000000100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1001000000100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1001000000100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1001000000100000100) && ({row_reg, col_reg}<19'b1001000000101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1001000000101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1001000000101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001000000110000000) && ({row_reg, col_reg}<19'b1001000000110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001000000110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1001000000110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1001000000110011010) && ({row_reg, col_reg}<19'b1001000010011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1001000010011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1001000010011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001000010011101010) && ({row_reg, col_reg}<19'b1001000010011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001000010011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1001000010011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001000010011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001000010011101111) && ({row_reg, col_reg}<19'b1001000010100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001000010100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1001000010100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1001000010100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1001000010100000100) && ({row_reg, col_reg}<19'b1001000010101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1001000010101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1001000010101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001000010110000000) && ({row_reg, col_reg}<19'b1001000010110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001000010110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1001000010110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1001000010110011010) && ({row_reg, col_reg}<19'b1001000100011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1001000100011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1001000100011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001000100011101010) && ({row_reg, col_reg}<19'b1001000100011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001000100011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1001000100011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001000100011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001000100011101111) && ({row_reg, col_reg}<19'b1001000100100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001000100100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1001000100100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1001000100100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1001000100100000100) && ({row_reg, col_reg}<19'b1001000100101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1001000100101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1001000100101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001000100110000000) && ({row_reg, col_reg}<19'b1001000100110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001000100110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1001000100110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1001000100110011010) && ({row_reg, col_reg}<19'b1001000110011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1001000110011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1001000110011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001000110011101010) && ({row_reg, col_reg}<19'b1001000110011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001000110011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1001000110011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001000110011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001000110011101111) && ({row_reg, col_reg}<19'b1001000110100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001000110100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1001000110100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1001000110100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1001000110100000100) && ({row_reg, col_reg}<19'b1001000110101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1001000110101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1001000110101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001000110110000000) && ({row_reg, col_reg}<19'b1001000110110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001000110110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1001000110110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1001000110110011010) && ({row_reg, col_reg}<19'b1001001000011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1001001000011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1001001000011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001001000011101010) && ({row_reg, col_reg}<19'b1001001000011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001001000011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1001001000011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001001000011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001001000011101111) && ({row_reg, col_reg}<19'b1001001000100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001001000100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1001001000100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1001001000100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1001001000100000100) && ({row_reg, col_reg}<19'b1001001000101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1001001000101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1001001000101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001001000110000000) && ({row_reg, col_reg}<19'b1001001000110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001001000110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1001001000110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1001001000110011010) && ({row_reg, col_reg}<19'b1001001010011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1001001010011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1001001010011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001001010011101010) && ({row_reg, col_reg}<19'b1001001010011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001001010011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1001001010011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001001010011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001001010011101111) && ({row_reg, col_reg}<19'b1001001010100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001001010100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1001001010100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1001001010100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1001001010100000100) && ({row_reg, col_reg}<19'b1001001010101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1001001010101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1001001010101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001001010110000000) && ({row_reg, col_reg}<19'b1001001010110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001001010110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1001001010110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1001001010110011010) && ({row_reg, col_reg}<19'b1001001100011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1001001100011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1001001100011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001001100011101010) && ({row_reg, col_reg}<19'b1001001100011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001001100011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1001001100011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001001100011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001001100011101111) && ({row_reg, col_reg}<19'b1001001100100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001001100100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1001001100100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1001001100100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1001001100100000100) && ({row_reg, col_reg}<19'b1001001100101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1001001100101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1001001100101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001001100110000000) && ({row_reg, col_reg}<19'b1001001100110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001001100110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1001001100110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1001001100110011010) && ({row_reg, col_reg}<19'b1001001110011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1001001110011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1001001110011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001001110011101010) && ({row_reg, col_reg}<19'b1001001110011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001001110011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1001001110011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001001110011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001001110011101111) && ({row_reg, col_reg}<19'b1001001110100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001001110100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1001001110100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1001001110100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1001001110100000100) && ({row_reg, col_reg}<19'b1001001110101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1001001110101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1001001110101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001001110110000000) && ({row_reg, col_reg}<19'b1001001110110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001001110110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1001001110110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1001001110110011010) && ({row_reg, col_reg}<19'b1001010000011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1001010000011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1001010000011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001010000011101010) && ({row_reg, col_reg}<19'b1001010000011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001010000011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1001010000011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001010000011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001010000011101111) && ({row_reg, col_reg}<19'b1001010000100000000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001010000100000000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1001010000100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001010000100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1001010000100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1001010000100000100) && ({row_reg, col_reg}<19'b1001010000101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1001010000101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1001010000101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001010000110000000) && ({row_reg, col_reg}<19'b1001010000110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001010000110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1001010000110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1001010000110011010) && ({row_reg, col_reg}<19'b1001010010011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1001010010011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1001010010011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001010010011101010) && ({row_reg, col_reg}<19'b1001010010011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001010010011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1001010010011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001010010011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001010010011101111) && ({row_reg, col_reg}<19'b1001010010100000000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001010010100000000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1001010010100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001010010100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1001010010100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1001010010100000100) && ({row_reg, col_reg}<19'b1001010010101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1001010010101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1001010010101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001010010110000000) && ({row_reg, col_reg}<19'b1001010010110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001010010110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1001010010110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1001010010110011010) && ({row_reg, col_reg}<19'b1001010100011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1001010100011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1001010100011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001010100011101010) && ({row_reg, col_reg}<19'b1001010100011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001010100011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1001010100011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001010100011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001010100011101111) && ({row_reg, col_reg}<19'b1001010100100000000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001010100100000000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1001010100100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001010100100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1001010100100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1001010100100000100) && ({row_reg, col_reg}<19'b1001010100101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1001010100101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1001010100101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001010100110000000) && ({row_reg, col_reg}<19'b1001010100110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001010100110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1001010100110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1001010100110011010) && ({row_reg, col_reg}<19'b1001010110011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1001010110011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1001010110011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001010110011101010) && ({row_reg, col_reg}<19'b1001010110011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001010110011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1001010110011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001010110011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001010110011101111) && ({row_reg, col_reg}<19'b1001010110100000000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001010110100000000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1001010110100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001010110100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1001010110100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1001010110100000100) && ({row_reg, col_reg}<19'b1001010110101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1001010110101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1001010110101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001010110110000000) && ({row_reg, col_reg}<19'b1001010110110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001010110110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1001010110110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1001010110110011010) && ({row_reg, col_reg}<19'b1001011000011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1001011000011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1001011000011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001011000011101010) && ({row_reg, col_reg}<19'b1001011000011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001011000011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1001011000011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001011000011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001011000011101111) && ({row_reg, col_reg}<19'b1001011000100000000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001011000100000000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1001011000100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001011000100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1001011000100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1001011000100000100) && ({row_reg, col_reg}<19'b1001011000101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1001011000101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1001011000101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001011000110000000) && ({row_reg, col_reg}<19'b1001011000110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001011000110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1001011000110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1001011000110011010) && ({row_reg, col_reg}<19'b1001011010011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1001011010011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1001011010011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001011010011101010) && ({row_reg, col_reg}<19'b1001011010011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001011010011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1001011010011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001011010011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001011010011101111) && ({row_reg, col_reg}<19'b1001011010100000000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001011010100000000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1001011010100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001011010100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1001011010100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1001011010100000100) && ({row_reg, col_reg}<19'b1001011010101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1001011010101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1001011010101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001011010110000000) && ({row_reg, col_reg}<19'b1001011010110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001011010110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1001011010110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1001011010110011010) && ({row_reg, col_reg}<19'b1001011100011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1001011100011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1001011100011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001011100011101010) && ({row_reg, col_reg}<19'b1001011100011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001011100011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1001011100011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001011100011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001011100011101111) && ({row_reg, col_reg}<19'b1001011100100000000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001011100100000000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1001011100100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001011100100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1001011100100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1001011100100000100) && ({row_reg, col_reg}<19'b1001011100101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1001011100101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1001011100101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001011100110000000) && ({row_reg, col_reg}<19'b1001011100110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001011100110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1001011100110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1001011100110011010) && ({row_reg, col_reg}<19'b1001011110011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1001011110011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1001011110011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001011110011101010) && ({row_reg, col_reg}<19'b1001011110011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001011110011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1001011110011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001011110011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001011110011101111) && ({row_reg, col_reg}<19'b1001011110100000000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001011110100000000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1001011110100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001011110100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1001011110100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1001011110100000100) && ({row_reg, col_reg}<19'b1001011110101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1001011110101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1001011110101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001011110110000000) && ({row_reg, col_reg}<19'b1001011110110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001011110110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1001011110110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1001011110110011010) && ({row_reg, col_reg}<19'b1001100000011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1001100000011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1001100000011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1001100000011101010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001100000011101011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001100000011101100) && ({row_reg, col_reg}<19'b1001100000100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001100000100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1001100000100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1001100000100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1001100000100000100) && ({row_reg, col_reg}<19'b1001100000101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1001100000101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1001100000101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001100000110000000) && ({row_reg, col_reg}<19'b1001100000110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001100000110011000)) color_data = 12'b101010101010;

		if(({row_reg, col_reg}>=19'b1001100000110011001) && ({row_reg, col_reg}<19'b1001100010011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1001100010011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1001100010011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001100010011101010) && ({row_reg, col_reg}<19'b1001100010100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001100010100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1001100010100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1001100010100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1001100010100000100) && ({row_reg, col_reg}<19'b1001100010101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1001100010101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1001100010101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001100010110000000) && ({row_reg, col_reg}<19'b1001100010110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001100010110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1001100010110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1001100010110011010) && ({row_reg, col_reg}<19'b1001100100001011001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1001100100001011001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=19'b1001100100001011010) && ({row_reg, col_reg}<19'b1001100100001011100)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1001100100001011100) && ({row_reg, col_reg}<19'b1001100100001011110)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=19'b1001100100001011110) && ({row_reg, col_reg}<19'b1001100100011101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1001100100011101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1001100100011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001100100011101010) && ({row_reg, col_reg}<19'b1001100100011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001100100011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1001100100011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001100100011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001100100011101111) && ({row_reg, col_reg}<19'b1001100100100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b1001100100100000001) && ({row_reg, col_reg}<19'b1001100100100000011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1001100100100000011)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=19'b1001100100100000100) && ({row_reg, col_reg}<19'b1001100100101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1001100100101111110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=19'b1001100100101111111) && ({row_reg, col_reg}<19'b1001100100110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001100100110011000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001100100110011001) && ({row_reg, col_reg}<19'b1001100101000100001)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=19'b1001100101000100001) && ({row_reg, col_reg}<19'b1001100101000100011)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1001100101000100011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1001100101000100100) && ({row_reg, col_reg}<19'b1001100101000100110)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1001100101000100110) && ({row_reg, col_reg}<19'b1001100110001010110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1001100110001010110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b1001100110001010111)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b1001100110001011000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1001100110001011001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1001100110001011010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=19'b1001100110001011011) && ({row_reg, col_reg}<19'b1001100110001011110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1001100110001011110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b1001100110001011111) && ({row_reg, col_reg}<19'b1001100110011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001100110011101001) && ({row_reg, col_reg}<19'b1001100110011101011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b1001100110011101011) && ({row_reg, col_reg}<19'b1001100110011101101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1001100110011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001100110011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001100110011101111) && ({row_reg, col_reg}<19'b1001100110100000000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b1001100110100000000) && ({row_reg, col_reg}<19'b1001100110100000010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1001100110100000010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b1001100110100000011) && ({row_reg, col_reg}<19'b1001100110110000000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001100110110000000) && ({row_reg, col_reg}<19'b1001100110110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b1001100110110011000) && ({row_reg, col_reg}<19'b1001100111000100011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001100111000100011) && ({row_reg, col_reg}<19'b1001100111000100101)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1001100111000100101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1001100111000100110)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1001100111000100111)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1001100111000101000) && ({row_reg, col_reg}<19'b1001101000001010101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1001101000001010101)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b1001101000001010110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1001101000001010111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1001101000001011000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001101000001011001) && ({row_reg, col_reg}<19'b1001101000001011011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b1001101000001011011) && ({row_reg, col_reg}<19'b1001101000001100000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001101000001100000) && ({row_reg, col_reg}<19'b1001101000011101001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001101000011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1001101000011101010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001101000011101011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001101000011101100) && ({row_reg, col_reg}<19'b1001101000011101110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b1001101000011101110) && ({row_reg, col_reg}<19'b1001101000011110000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001101000011110000) && ({row_reg, col_reg}<19'b1001101000100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001101000100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1001101000100000010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001101000100000011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1001101000100000100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001101000100000101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001101000100000110) && ({row_reg, col_reg}<19'b1001101000101111000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b1001101000101111000) && ({row_reg, col_reg}<19'b1001101000101111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001101000101111010) && ({row_reg, col_reg}<19'b1001101000101111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001101000101111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001101000101111101) && ({row_reg, col_reg}<19'b1001101000110011101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001101000110011101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001101000110011110) && ({row_reg, col_reg}<19'b1001101001000100000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001101001000100000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001101001000100001) && ({row_reg, col_reg}<19'b1001101001000100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001101001000100110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1001101001000100111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1001101001000101000)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b1001101001000101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1001101001000101010) && ({row_reg, col_reg}<19'b1001101010001010100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1001101010001010100)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b1001101010001010101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1001101010001010110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001101010001010111) && ({row_reg, col_reg}<19'b1001101010001011011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b1001101010001011011) && ({row_reg, col_reg}<19'b1001101010001011101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001101010001011101) && ({row_reg, col_reg}<19'b1001101010001100000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b1001101010001100000) && ({row_reg, col_reg}<19'b1001101010011101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1001101010011101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001101010011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1001101010011101010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001101010011101011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1001101010011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001101010011101101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001101010011101110) && ({row_reg, col_reg}<19'b1001101010100000010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001101010100000010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001101010100000011) && ({row_reg, col_reg}<19'b1001101010100001000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b1001101010100001000) && ({row_reg, col_reg}<19'b1001101010101111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001101010101111001) && ({row_reg, col_reg}<19'b1001101010101111011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b1001101010101111011) && ({row_reg, col_reg}<19'b1001101010101111101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001101010101111101) && ({row_reg, col_reg}<19'b1001101010110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b1001101010110011000) && ({row_reg, col_reg}<19'b1001101010110011110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1001101010110011110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b1001101010110011111) && ({row_reg, col_reg}<19'b1001101011000100000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001101011000100000) && ({row_reg, col_reg}<19'b1001101011000100111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001101011000100111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1001101011000101000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1001101011000101001)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1001101011000101010)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1001101011000101011) && ({row_reg, col_reg}<19'b1001101100001010011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1001101100001010011)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1001101100001010100)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=19'b1001101100001010101) && ({row_reg, col_reg}<19'b1001101100001010111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b1001101100001010111) && ({row_reg, col_reg}<19'b1001101100001011011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001101100001011011) && ({row_reg, col_reg}<19'b1001101100001011110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b1001101100001011110) && ({row_reg, col_reg}<19'b1001101100001100000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001101100001100000) && ({row_reg, col_reg}<19'b1001101100011101011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001101100011101011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1001101100011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001101100011101101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001101100011101110) && ({row_reg, col_reg}<19'b1001101100100000000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b1001101100100000000) && ({row_reg, col_reg}<19'b1001101100100000011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001101100100000011) && ({row_reg, col_reg}<19'b1001101100100000101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b1001101100100000101) && ({row_reg, col_reg}<19'b1001101100100001000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001101100100001000) && ({row_reg, col_reg}<19'b1001101100101111011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001101100101111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1001101100101111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b1001101100101111101) && ({row_reg, col_reg}<19'b1001101100110000000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001101100110000000) && ({row_reg, col_reg}<19'b1001101100110011110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b1001101100110011110) && ({row_reg, col_reg}<19'b1001101100110100000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001101100110100000) && ({row_reg, col_reg}<19'b1001101101000100000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b1001101101000100000) && ({row_reg, col_reg}<19'b1001101101000100011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001101101000100011) && ({row_reg, col_reg}<19'b1001101101000100101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b1001101101000100101) && ({row_reg, col_reg}<19'b1001101101000100111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001101101000100111) && ({row_reg, col_reg}<19'b1001101101000101001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001101101000101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1001101101000101010)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1001101101000101011)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1001101101000101100) && ({row_reg, col_reg}<19'b1001101110001010010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1001101110001010010)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b1001101110001010011)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=19'b1001101110001010100) && ({row_reg, col_reg}<19'b1001101110001010110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001101110001010110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001101110001010111) && ({row_reg, col_reg}<19'b1001101110001011010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001101110001011010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001101110001011011) && ({row_reg, col_reg}<19'b1001101110001011101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b1001101110001011101) && ({row_reg, col_reg}<19'b1001101110001011111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001101110001011111) && ({row_reg, col_reg}<19'b1001101110011101011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001101110011101011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1001101110011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001101110011101101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1001101110011101110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001101110011101111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001101110011110000) && ({row_reg, col_reg}<19'b1001101110100000000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001101110100000000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001101110100000001) && ({row_reg, col_reg}<19'b1001101110100000100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b1001101110100000100) && ({row_reg, col_reg}<19'b1001101110100000110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001101110100000110) && ({row_reg, col_reg}<19'b1001101110101111000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b1001101110101111000) && ({row_reg, col_reg}<19'b1001101110101111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1001101110101111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001101110101111101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001101110101111110) && ({row_reg, col_reg}<19'b1001101110110011001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001101110110011001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001101110110011010) && ({row_reg, col_reg}<19'b1001101110110011100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b1001101110110011100) && ({row_reg, col_reg}<19'b1001101110110011111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001101110110011111) && ({row_reg, col_reg}<19'b1001101111000101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001101111000101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1001101111000101001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001101111000101010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1001101111000101011)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=19'b1001101111000101100) && ({row_reg, col_reg}<19'b1001110000001010001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1001110000001010001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b1001110000001010010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1001110000001010011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001110000001010100) && ({row_reg, col_reg}<19'b1001110000001010110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001110000001010110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001110000001010111) && ({row_reg, col_reg}<19'b1001110001000101001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b1001110001000101001) && ({row_reg, col_reg}<19'b1001110001000101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1001110001000101100)) color_data = 12'b110111011101;

		if(({row_reg, col_reg}>=19'b1001110001000101101) && ({row_reg, col_reg}<19'b1001110010001010001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1001110010001010001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1001110010001010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1001110010001010011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001110010001010100) && ({row_reg, col_reg}<19'b1001110010001010110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001110010001010110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001110010001010111) && ({row_reg, col_reg}<19'b1001110011000101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001110011000101100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1001110011000101101)) color_data = 12'b110111011101;

		if(({row_reg, col_reg}>=19'b1001110011000101110) && ({row_reg, col_reg}<19'b1001110100001010000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1001110100001010000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b1001110100001010001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=19'b1001110100001010010) && ({row_reg, col_reg}<19'b1001110100001010100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b1001110100001010100) && ({row_reg, col_reg}<19'b1001110100001010111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001110100001010111) && ({row_reg, col_reg}<19'b1001110101000101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001110101000101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001110101000101001) && ({row_reg, col_reg}<19'b1001110101000101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001110101000101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1001110101000101101)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=19'b1001110101000101110) && ({row_reg, col_reg}<19'b1001110110001010000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1001110110001010000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1001110110001010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1001110110001010010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001110110001010011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1001110110001010100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b1001110110001010101) && ({row_reg, col_reg}<19'b1001110110001010111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001110110001010111) && ({row_reg, col_reg}<19'b1001110111000101001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b1001110111000101001) && ({row_reg, col_reg}<19'b1001110111000101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1001110111000101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001110111000101101)) color_data = 12'b101110111011;

		if(({row_reg, col_reg}>=19'b1001110111000101110) && ({row_reg, col_reg}<19'b1001111000001010000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1001111000001010000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1001111000001010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1001111000001010010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001111000001010011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1001111000001010100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001111000001010101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001111000001010110) && ({row_reg, col_reg}<19'b1001111001000101001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b1001111001000101001) && ({row_reg, col_reg}<19'b1001111001000101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1001111001000101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001111001000101101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1001111001000101110)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1001111001000101111) && ({row_reg, col_reg}<19'b1001111010001010000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1001111010001010000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1001111010001010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1001111010001010010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001111010001010011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001111010001010100) && ({row_reg, col_reg}<19'b1001111010001010111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001111010001010111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001111010001011000) && ({row_reg, col_reg}<19'b1001111011000101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b1001111011000101000) && ({row_reg, col_reg}<19'b1001111011000101010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001111011000101010) && ({row_reg, col_reg}<19'b1001111011000101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001111011000101101)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1001111011000101110)) color_data = 12'b110111011101;

		if(({row_reg, col_reg}>=19'b1001111011000101111) && ({row_reg, col_reg}<19'b1001111100001010000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1001111100001010000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1001111100001010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001111100001010010) && ({row_reg, col_reg}<19'b1001111100001010100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b1001111100001010100) && ({row_reg, col_reg}<19'b1001111100001010110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1001111100001010110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001111100001010111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001111100001011000) && ({row_reg, col_reg}<19'b1001111101000101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001111101000101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1001111101000101001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001111101000101010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001111101000101011) && ({row_reg, col_reg}<19'b1001111101000101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001111101000101101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1001111101000101110)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=19'b1001111101000101111) && ({row_reg, col_reg}<19'b1001111110001010000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=19'b1001111110001010000) && ({row_reg, col_reg}<19'b1001111110001010010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001111110001010010) && ({row_reg, col_reg}<19'b1001111110001010100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b1001111110001010100) && ({row_reg, col_reg}<19'b1001111110001010110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001111110001010110) && ({row_reg, col_reg}<19'b1001111111000101010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001111111000101010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001111111000101011) && ({row_reg, col_reg}<19'b1001111111000101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001111111000101101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1001111111000101110)) color_data = 12'b101110111011;

		if(({row_reg, col_reg}>=19'b1001111111000101111) && ({row_reg, col_reg}<19'b1010000000001010000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=19'b1010000000001010000) && ({row_reg, col_reg}<19'b1010000000001010010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1010000000001010010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010000000001010011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1010000000001010100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b1010000000001010101) && ({row_reg, col_reg}<19'b1010000000001010111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010000000001010111) && ({row_reg, col_reg}<19'b1010000001000101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010000001000101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1010000001000101001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010000001000101010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010000001000101011) && ({row_reg, col_reg}<19'b1010000001000101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010000001000101101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1010000001000101110)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=19'b1010000001000101111) && ({row_reg, col_reg}<19'b1010000010001010000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1010000010001010000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1010000010001010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010000010001010010) && ({row_reg, col_reg}<19'b1010000010001010101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b1010000010001010101) && ({row_reg, col_reg}<19'b1010000010001011000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010000010001011000) && ({row_reg, col_reg}<19'b1010000011000101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010000011000101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1010000011000101001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010000011000101010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1010000011000101011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b1010000011000101100) && ({row_reg, col_reg}<19'b1010000011000101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1010000011000101110)) color_data = 12'b110111011101;

		if(({row_reg, col_reg}>=19'b1010000011000101111) && ({row_reg, col_reg}<19'b1010000100001010000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1010000100001010000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=19'b1010000100001010001) && ({row_reg, col_reg}<19'b1010000100001010011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010000100001010011) && ({row_reg, col_reg}<19'b1010000100001010101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010000100001010101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1010000100001010110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010000100001010111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010000100001011000) && ({row_reg, col_reg}<19'b1010000101000101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b1010000101000101000) && ({row_reg, col_reg}<19'b1010000101000101010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010000101000101010) && ({row_reg, col_reg}<19'b1010000101000101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010000101000101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1010000101000101101)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1010000101000101110)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1010000101000101111) && ({row_reg, col_reg}<19'b1010000110001010000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1010000110001010000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=19'b1010000110001010001) && ({row_reg, col_reg}<19'b1010000110001010101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010000110001010101) && ({row_reg, col_reg}<19'b1010000110001010111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010000110001010111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010000110001011000) && ({row_reg, col_reg}<19'b1010000111000101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010000111000101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1010000111000101101)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1010000111000101110)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1010000111000101111) && ({row_reg, col_reg}<19'b1010001000001010000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1010001000001010000)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b1010001000001010001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1010001000001010010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b1010001000001010011) && ({row_reg, col_reg}<19'b1010001000001010110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1010001000001010110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010001000001010111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010001000001011000) && ({row_reg, col_reg}<19'b1010001001000101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010001001000101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1010001001000101101)) color_data = 12'b101110111011;

		if(({row_reg, col_reg}>=19'b1010001001000101110) && ({row_reg, col_reg}<19'b1010001010001010000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1010001010001010000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b1010001010001010001)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1010001010001010010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010001010001010011) && ({row_reg, col_reg}<19'b1010001010001010101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b1010001010001010101) && ({row_reg, col_reg}<19'b1010001010001010111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010001010001010111) && ({row_reg, col_reg}<19'b1010001011000101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010001011000101100)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1010001011000101101)) color_data = 12'b110111011101;

		if(({row_reg, col_reg}>=19'b1010001011000101110) && ({row_reg, col_reg}<19'b1010001100001010001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1010001100001010001)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b1010001100001010010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1010001100001010011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010001100001010100) && ({row_reg, col_reg}<19'b1010001101000101010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010001101000101010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1010001101000101011)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1010001101000101100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=19'b1010001101000101101) && ({row_reg, col_reg}<19'b1010001110001010010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1010001110001010010)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1010001110001010011)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1010001110001010100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010001110001010101) && ({row_reg, col_reg}<19'b1010001111000101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010001111000101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1010001111000101001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010001111000101010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1010001111000101011)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1010001111000101100)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1010001111000101101) && ({row_reg, col_reg}<19'b1010010000001010011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1010010000001010011)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1010010000001010100)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1010010000001010101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b1010010000001010110) && ({row_reg, col_reg}<19'b1010010000001100000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010010000001100000) && ({row_reg, col_reg}<19'b1010010000011101010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b1010010000011101010) && ({row_reg, col_reg}<19'b1010010000011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1010010000011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b1010010000011101101) && ({row_reg, col_reg}<19'b1010010000011101111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010010000011101111) && ({row_reg, col_reg}<19'b1010010000100000000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010010000100000000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1010010000100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010010000100000010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010010000100000011) && ({row_reg, col_reg}<19'b1010010000100000101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b1010010000100000101) && ({row_reg, col_reg}<19'b1010010000100000111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010010000100000111) && ({row_reg, col_reg}<19'b1010010000101111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010010000101111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010010000101111011) && ({row_reg, col_reg}<19'b1010010000110011001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010010000110011001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010010000110011010) && ({row_reg, col_reg}<19'b1010010000110011100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010010000110011100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010010000110011101) && ({row_reg, col_reg}<19'b1010010000110011111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010010000110011111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010010000110100000) && ({row_reg, col_reg}<19'b1010010001000100001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b1010010001000100001) && ({row_reg, col_reg}<19'b1010010001000100011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1010010001000100011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b1010010001000100100) && ({row_reg, col_reg}<19'b1010010001000100110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010010001000100110) && ({row_reg, col_reg}<19'b1010010001000101001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010010001000101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1010010001000101010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1010010001000101011)) color_data = 12'b110111011101;

		if(({row_reg, col_reg}>=19'b1010010001000101100) && ({row_reg, col_reg}<19'b1010010010001010011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1010010010001010011)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b1010010010001010100)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1010010010001010101)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1010010010001010110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010010010001010111) && ({row_reg, col_reg}<19'b1010010010001011100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010010010001011100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010010010001011101) && ({row_reg, col_reg}<19'b1010010010011101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010010010011101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010010010011101001) && ({row_reg, col_reg}<19'b1010010010011101011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010010010011101011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1010010010011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010010010011101101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010010010011101110) && ({row_reg, col_reg}<19'b1010010010100000010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b1010010010100000010) && ({row_reg, col_reg}<19'b1010010010100000101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010010010100000101) && ({row_reg, col_reg}<19'b1010010010100000111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010010010100000111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010010010100001000) && ({row_reg, col_reg}<19'b1010010010101111000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010010010101111000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010010010101111001) && ({row_reg, col_reg}<19'b1010010010101111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b1010010010101111101) && ({row_reg, col_reg}<19'b1010010010110000000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010010010110000000) && ({row_reg, col_reg}<19'b1010010010110011001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b1010010010110011001) && ({row_reg, col_reg}<19'b1010010010110011101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010010010110011101) && ({row_reg, col_reg}<19'b1010010011000100000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010010011000100000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010010011000100001) && ({row_reg, col_reg}<19'b1010010011000100011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b1010010011000100011) && ({row_reg, col_reg}<19'b1010010011000100101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010010011000100101) && ({row_reg, col_reg}<19'b1010010011000100111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b1010010011000100111) && ({row_reg, col_reg}<19'b1010010011000101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1010010011000101001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1010010011000101010)) color_data = 12'b110111011101;

		if(({row_reg, col_reg}>=19'b1010010011000101011) && ({row_reg, col_reg}<19'b1010010100001010100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1010010100001010100)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b1010010100001010101)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b1010010100001010110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=19'b1010010100001010111) && ({row_reg, col_reg}<19'b1010010100001011010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010010100001011010) && ({row_reg, col_reg}<19'b1010010100001011100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b1010010100001011100) && ({row_reg, col_reg}<19'b1010010100011100000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010010100011100000) && ({row_reg, col_reg}<19'b1010010100011101010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010010100011101010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010010100011101011) && ({row_reg, col_reg}<19'b1010010100100000000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b1010010100100000000) && ({row_reg, col_reg}<19'b1010010100100000100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010010100100000100) && ({row_reg, col_reg}<19'b1010010100100001000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b1010010100100001000) && ({row_reg, col_reg}<19'b1010010100101111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010010100101111001) && ({row_reg, col_reg}<19'b1010010100101111011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b1010010100101111011) && ({row_reg, col_reg}<19'b1010010100101111101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010010100101111101) && ({row_reg, col_reg}<19'b1010010100110011001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b1010010100110011001) && ({row_reg, col_reg}<19'b1010010100110011011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1010010100110011011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010010100110011100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1010010100110011101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010010100110011110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1010010100110011111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b1010010100110100000) && ({row_reg, col_reg}<19'b1010010101000100000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010010101000100000) && ({row_reg, col_reg}<19'b1010010101000100011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010010101000100011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010010101000100100) && ({row_reg, col_reg}<19'b1010010101000100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010010101000100110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1010010101000100111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1010010101000101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1010010101000101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1010010101000101010) && ({row_reg, col_reg}<19'b1010010110001010110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1010010110001010110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b1010010110001010111)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=19'b1010010110001011000) && ({row_reg, col_reg}<19'b1010010110001011010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=19'b1010010110001011010) && ({row_reg, col_reg}<19'b1010010110001011101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010010110001011101) && ({row_reg, col_reg}<19'b1010010110001011111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010010110001011111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010010110001100000) && ({row_reg, col_reg}<19'b1010010110011101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010010110011101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1010010110011101001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010010110011101010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010010110011101011) && ({row_reg, col_reg}<19'b1010010110011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b1010010110011101101) && ({row_reg, col_reg}<19'b1010010110011101111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010010110011101111) && ({row_reg, col_reg}<19'b1010010110100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010010110100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1010010110100000010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010010110100000011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1010010110100000100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b1010010110100000101) && ({row_reg, col_reg}<19'b1010010110100000111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010010110100000111) && ({row_reg, col_reg}<19'b1010010110101111000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010010110101111000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010010110101111001) && ({row_reg, col_reg}<19'b1010010110101111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010010110101111101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1010010110101111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010010110101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010010110110000000) && ({row_reg, col_reg}<19'b1010010110110011001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010010110110011001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010010110110011010) && ({row_reg, col_reg}<19'b1010010110110011110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010010110110011110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010010110110011111) && ({row_reg, col_reg}<19'b1010010111000100000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b1010010111000100000) && ({row_reg, col_reg}<19'b1010010111000100101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1010010111000100101)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1010010111000100110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1010010111000100111)) color_data = 12'b110111011101;

		if(({row_reg, col_reg}>=19'b1010010111000101000) && ({row_reg, col_reg}<19'b1010011000001011000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1010011000001011000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b1010011000001011001)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b1010011000001011010)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1010011000001011011)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=19'b1010011000001011100) && ({row_reg, col_reg}<19'b1010011000001011110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1010011000001011110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=19'b1010011000001011111) && ({row_reg, col_reg}<19'b1010011000011101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1010011000011101000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=19'b1010011000011101001) && ({row_reg, col_reg}<19'b1010011000011101011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010011000011101011) && ({row_reg, col_reg}<19'b1010011000011101111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010011000011101111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010011000011110000) && ({row_reg, col_reg}<19'b1010011000100000010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010011000100000010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1010011000100000011)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=19'b1010011000100000100) && ({row_reg, col_reg}<19'b1010011000100000111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1010011000100000111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=19'b1010011000100001000) && ({row_reg, col_reg}<19'b1010011000101111000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=19'b1010011000101111000) && ({row_reg, col_reg}<19'b1010011000101111010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1010011000101111010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=19'b1010011000101111011) && ({row_reg, col_reg}<19'b1010011000101111101)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1010011000101111101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=19'b1010011000101111110) && ({row_reg, col_reg}<19'b1010011000110000000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010011000110000000) && ({row_reg, col_reg}<19'b1010011000110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010011000110011000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1010011000110011001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1010011000110011010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1010011000110011011)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1010011000110011100)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=19'b1010011000110011101) && ({row_reg, col_reg}<19'b1010011000110011111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1010011000110011111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=19'b1010011000110100000) && ({row_reg, col_reg}<19'b1010011001000100000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1010011001000100000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1010011001000100001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1010011001000100010)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1010011001000100011)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=19'b1010011001000100100) && ({row_reg, col_reg}<19'b1010011001000100110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b1010011001000100110)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1010011001000100111) && ({row_reg, col_reg}<19'b1010011010001011110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=19'b1010011010001011110) && ({row_reg, col_reg}<19'b1010011010011101000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b1010011010011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1010011010011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010011010011101010) && ({row_reg, col_reg}<19'b1010011010011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010011010011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010011010011101101) && ({row_reg, col_reg}<19'b1010011010011101111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010011010011101111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010011010011110000) && ({row_reg, col_reg}<19'b1010011010100000000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b1010011010100000000) && ({row_reg, col_reg}<19'b1010011010100000010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1010011010100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1010011010100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1010011010100000100) && ({row_reg, col_reg}<19'b1010011010101111110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b1010011010101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1010011010101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010011010110000000) && ({row_reg, col_reg}<19'b1010011010110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010011010110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1010011010110011001)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b1010011010110011010)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b1010011010110011011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=19'b1010011010110011100) && ({row_reg, col_reg}<19'b1010011011000100000)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1010011011000100000) && ({row_reg, col_reg}<19'b1010011100011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1010011100011101000)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b1010011100011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010011100011101010) && ({row_reg, col_reg}<19'b1010011100011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010011100011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010011100011101101) && ({row_reg, col_reg}<19'b1010011100100000010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010011100100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1010011100100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1010011100100000100) && ({row_reg, col_reg}<19'b1010011100101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1010011100101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1010011100101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010011100110000000) && ({row_reg, col_reg}<19'b1010011100110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010011100110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1010011100110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1010011100110011010) && ({row_reg, col_reg}<19'b1010011110011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1010011110011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=19'b1010011110011101001) && ({row_reg, col_reg}<19'b1010011110011101011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010011110011101011) && ({row_reg, col_reg}<19'b1010011110011101110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010011110011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010011110011101111) && ({row_reg, col_reg}<19'b1010011110100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010011110100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1010011110100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1010011110100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1010011110100000100) && ({row_reg, col_reg}<19'b1010011110101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1010011110101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1010011110101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010011110110000000) && ({row_reg, col_reg}<19'b1010011110110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010011110110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1010011110110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1010011110110011010) && ({row_reg, col_reg}<19'b1010100000011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1010100000011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1010100000011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010100000011101010) && ({row_reg, col_reg}<19'b1010100000011101110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010100000011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010100000011101111) && ({row_reg, col_reg}<19'b1010100000100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010100000100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1010100000100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1010100000100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1010100000100000100) && ({row_reg, col_reg}<19'b1010100000101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1010100000101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1010100000101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010100000110000000) && ({row_reg, col_reg}<19'b1010100000110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010100000110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1010100000110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1010100000110011010) && ({row_reg, col_reg}<19'b1010100010011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1010100010011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1010100010011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010100010011101010) && ({row_reg, col_reg}<19'b1010100010011101110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010100010011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010100010011101111) && ({row_reg, col_reg}<19'b1010100010100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010100010100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1010100010100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1010100010100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1010100010100000100) && ({row_reg, col_reg}<19'b1010100010101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1010100010101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1010100010101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010100010110000000) && ({row_reg, col_reg}<19'b1010100010110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010100010110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1010100010110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1010100010110011010) && ({row_reg, col_reg}<19'b1010100100011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1010100100011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1010100100011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010100100011101010) && ({row_reg, col_reg}<19'b1010100100011101110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010100100011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010100100011101111) && ({row_reg, col_reg}<19'b1010100100100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010100100100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1010100100100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1010100100100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1010100100100000100) && ({row_reg, col_reg}<19'b1010100100101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1010100100101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1010100100101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010100100110000000) && ({row_reg, col_reg}<19'b1010100100110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010100100110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1010100100110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1010100100110011010) && ({row_reg, col_reg}<19'b1010100110011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1010100110011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1010100110011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010100110011101010) && ({row_reg, col_reg}<19'b1010100110011101110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010100110011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010100110011101111) && ({row_reg, col_reg}<19'b1010100110100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010100110100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1010100110100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1010100110100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1010100110100000100) && ({row_reg, col_reg}<19'b1010100110101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1010100110101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1010100110101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010100110110000000) && ({row_reg, col_reg}<19'b1010100110110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010100110110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1010100110110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1010100110110011010) && ({row_reg, col_reg}<19'b1010101000011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1010101000011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1010101000011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010101000011101010) && ({row_reg, col_reg}<19'b1010101000011101110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010101000011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010101000011101111) && ({row_reg, col_reg}<19'b1010101000100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010101000100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1010101000100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1010101000100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1010101000100000100) && ({row_reg, col_reg}<19'b1010101000101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1010101000101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1010101000101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010101000110000000) && ({row_reg, col_reg}<19'b1010101000110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010101000110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1010101000110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1010101000110011010) && ({row_reg, col_reg}<19'b1010101010011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1010101010011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1010101010011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010101010011101010) && ({row_reg, col_reg}<19'b1010101010011101110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010101010011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010101010011101111) && ({row_reg, col_reg}<19'b1010101010100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010101010100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1010101010100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1010101010100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1010101010100000100) && ({row_reg, col_reg}<19'b1010101010101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1010101010101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1010101010101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010101010110000000) && ({row_reg, col_reg}<19'b1010101010110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010101010110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1010101010110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1010101010110011010) && ({row_reg, col_reg}<19'b1010101100011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1010101100011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1010101100011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010101100011101010) && ({row_reg, col_reg}<19'b1010101100011101110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010101100011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010101100011101111) && ({row_reg, col_reg}<19'b1010101100100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010101100100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1010101100100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1010101100100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1010101100100000100) && ({row_reg, col_reg}<19'b1010101100101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1010101100101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1010101100101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010101100110000000) && ({row_reg, col_reg}<19'b1010101100110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010101100110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1010101100110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1010101100110011010) && ({row_reg, col_reg}<19'b1010101110011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1010101110011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1010101110011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010101110011101010) && ({row_reg, col_reg}<19'b1010101110011101110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010101110011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010101110011101111) && ({row_reg, col_reg}<19'b1010101110100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010101110100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1010101110100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1010101110100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1010101110100000100) && ({row_reg, col_reg}<19'b1010101110101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1010101110101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1010101110101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010101110110000000) && ({row_reg, col_reg}<19'b1010101110110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010101110110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1010101110110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1010101110110011010) && ({row_reg, col_reg}<19'b1010110000011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1010110000011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1010110000011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010110000011101010) && ({row_reg, col_reg}<19'b1010110000011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010110000011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1010110000011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010110000011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010110000011101111) && ({row_reg, col_reg}<19'b1010110000100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010110000100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1010110000100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1010110000100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1010110000100000100) && ({row_reg, col_reg}<19'b1010110000101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1010110000101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1010110000101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010110000110000000) && ({row_reg, col_reg}<19'b1010110000110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010110000110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1010110000110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1010110000110011010) && ({row_reg, col_reg}<19'b1010110010011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1010110010011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1010110010011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010110010011101010) && ({row_reg, col_reg}<19'b1010110010011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010110010011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1010110010011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010110010011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010110010011101111) && ({row_reg, col_reg}<19'b1010110010100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010110010100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1010110010100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1010110010100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1010110010100000100) && ({row_reg, col_reg}<19'b1010110010101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1010110010101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1010110010101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010110010110000000) && ({row_reg, col_reg}<19'b1010110010110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010110010110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1010110010110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1010110010110011010) && ({row_reg, col_reg}<19'b1010110100011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1010110100011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1010110100011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010110100011101010) && ({row_reg, col_reg}<19'b1010110100011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010110100011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1010110100011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010110100011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010110100011101111) && ({row_reg, col_reg}<19'b1010110100100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010110100100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1010110100100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1010110100100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1010110100100000100) && ({row_reg, col_reg}<19'b1010110100101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1010110100101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1010110100101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010110100110000000) && ({row_reg, col_reg}<19'b1010110100110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010110100110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1010110100110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1010110100110011010) && ({row_reg, col_reg}<19'b1010110110011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1010110110011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1010110110011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010110110011101010) && ({row_reg, col_reg}<19'b1010110110011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010110110011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1010110110011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010110110011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010110110011101111) && ({row_reg, col_reg}<19'b1010110110100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010110110100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1010110110100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1010110110100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1010110110100000100) && ({row_reg, col_reg}<19'b1010110110101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1010110110101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1010110110101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010110110110000000) && ({row_reg, col_reg}<19'b1010110110110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010110110110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1010110110110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1010110110110011010) && ({row_reg, col_reg}<19'b1010111000011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1010111000011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1010111000011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010111000011101010) && ({row_reg, col_reg}<19'b1010111000011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010111000011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1010111000011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010111000011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010111000011101111) && ({row_reg, col_reg}<19'b1010111000100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010111000100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1010111000100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1010111000100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1010111000100000100) && ({row_reg, col_reg}<19'b1010111000101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1010111000101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1010111000101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010111000110000000) && ({row_reg, col_reg}<19'b1010111000110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010111000110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1010111000110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1010111000110011010) && ({row_reg, col_reg}<19'b1010111010011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1010111010011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1010111010011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010111010011101010) && ({row_reg, col_reg}<19'b1010111010011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010111010011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1010111010011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010111010011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010111010011101111) && ({row_reg, col_reg}<19'b1010111010100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010111010100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1010111010100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1010111010100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1010111010100000100) && ({row_reg, col_reg}<19'b1010111010101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1010111010101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1010111010101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010111010110000000) && ({row_reg, col_reg}<19'b1010111010110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010111010110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1010111010110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1010111010110011010) && ({row_reg, col_reg}<19'b1010111100011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1010111100011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1010111100011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010111100011101010) && ({row_reg, col_reg}<19'b1010111100011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010111100011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1010111100011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010111100011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010111100011101111) && ({row_reg, col_reg}<19'b1010111100100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010111100100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1010111100100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1010111100100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1010111100100000100) && ({row_reg, col_reg}<19'b1010111100101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1010111100101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1010111100101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010111100110000000) && ({row_reg, col_reg}<19'b1010111100110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010111100110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1010111100110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1010111100110011010) && ({row_reg, col_reg}<19'b1010111110011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1010111110011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1010111110011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010111110011101010) && ({row_reg, col_reg}<19'b1010111110011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010111110011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1010111110011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010111110011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010111110011101111) && ({row_reg, col_reg}<19'b1010111110100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010111110100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1010111110100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1010111110100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1010111110100000100) && ({row_reg, col_reg}<19'b1010111110101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1010111110101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1010111110101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010111110110000000) && ({row_reg, col_reg}<19'b1010111110110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010111110110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1010111110110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1010111110110011010) && ({row_reg, col_reg}<19'b1011000000011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1011000000011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1011000000011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1011000000011101010) && ({row_reg, col_reg}<19'b1011000000011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011000000011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1011000000011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011000000011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1011000000011101111) && ({row_reg, col_reg}<19'b1011000000100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011000000100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1011000000100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1011000000100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1011000000100000100) && ({row_reg, col_reg}<19'b1011000000101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1011000000101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1011000000101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1011000000110000000) && ({row_reg, col_reg}<19'b1011000000110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011000000110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1011000000110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1011000000110011010) && ({row_reg, col_reg}<19'b1011000010011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1011000010011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1011000010011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1011000010011101010) && ({row_reg, col_reg}<19'b1011000010011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011000010011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1011000010011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011000010011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1011000010011101111) && ({row_reg, col_reg}<19'b1011000010100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011000010100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1011000010100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1011000010100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1011000010100000100) && ({row_reg, col_reg}<19'b1011000010101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1011000010101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1011000010101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1011000010110000000) && ({row_reg, col_reg}<19'b1011000010110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011000010110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1011000010110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1011000010110011010) && ({row_reg, col_reg}<19'b1011000100011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1011000100011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1011000100011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1011000100011101010) && ({row_reg, col_reg}<19'b1011000100011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011000100011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1011000100011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011000100011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1011000100011101111) && ({row_reg, col_reg}<19'b1011000100100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011000100100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1011000100100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1011000100100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1011000100100000100) && ({row_reg, col_reg}<19'b1011000100101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1011000100101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1011000100101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1011000100110000000) && ({row_reg, col_reg}<19'b1011000100110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011000100110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1011000100110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1011000100110011010) && ({row_reg, col_reg}<19'b1011000110011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1011000110011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1011000110011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1011000110011101010) && ({row_reg, col_reg}<19'b1011000110011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011000110011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1011000110011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011000110011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1011000110011101111) && ({row_reg, col_reg}<19'b1011000110100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011000110100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1011000110100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1011000110100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1011000110100000100) && ({row_reg, col_reg}<19'b1011000110101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1011000110101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1011000110101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1011000110110000000) && ({row_reg, col_reg}<19'b1011000110110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011000110110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1011000110110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1011000110110011010) && ({row_reg, col_reg}<19'b1011001000011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1011001000011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1011001000011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1011001000011101010) && ({row_reg, col_reg}<19'b1011001000011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011001000011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1011001000011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011001000011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1011001000011101111) && ({row_reg, col_reg}<19'b1011001000100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011001000100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1011001000100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1011001000100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1011001000100000100) && ({row_reg, col_reg}<19'b1011001000101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1011001000101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1011001000101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1011001000110000000) && ({row_reg, col_reg}<19'b1011001000110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011001000110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1011001000110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1011001000110011010) && ({row_reg, col_reg}<19'b1011001010011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1011001010011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1011001010011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1011001010011101010) && ({row_reg, col_reg}<19'b1011001010011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011001010011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1011001010011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011001010011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1011001010011101111) && ({row_reg, col_reg}<19'b1011001010100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011001010100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1011001010100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1011001010100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1011001010100000100) && ({row_reg, col_reg}<19'b1011001010101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1011001010101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1011001010101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1011001010110000000) && ({row_reg, col_reg}<19'b1011001010110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011001010110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1011001010110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1011001010110011010) && ({row_reg, col_reg}<19'b1011001100011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1011001100011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1011001100011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1011001100011101010) && ({row_reg, col_reg}<19'b1011001100011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011001100011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1011001100011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011001100011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1011001100011101111) && ({row_reg, col_reg}<19'b1011001100100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011001100100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1011001100100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1011001100100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1011001100100000100) && ({row_reg, col_reg}<19'b1011001100101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1011001100101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1011001100101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1011001100110000000) && ({row_reg, col_reg}<19'b1011001100110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011001100110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1011001100110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1011001100110011010) && ({row_reg, col_reg}<19'b1011001110011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1011001110011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1011001110011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1011001110011101010) && ({row_reg, col_reg}<19'b1011001110011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011001110011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1011001110011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011001110011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1011001110011101111) && ({row_reg, col_reg}<19'b1011001110100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011001110100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1011001110100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1011001110100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1011001110100000100) && ({row_reg, col_reg}<19'b1011001110101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1011001110101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1011001110101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1011001110110000000) && ({row_reg, col_reg}<19'b1011001110110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011001110110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1011001110110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1011001110110011010) && ({row_reg, col_reg}<19'b1011010000011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1011010000011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1011010000011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1011010000011101010) && ({row_reg, col_reg}<19'b1011010000011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011010000011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1011010000011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011010000011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1011010000011101111) && ({row_reg, col_reg}<19'b1011010000100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011010000100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1011010000100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1011010000100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1011010000100000100) && ({row_reg, col_reg}<19'b1011010000101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1011010000101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1011010000101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1011010000110000000) && ({row_reg, col_reg}<19'b1011010000110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011010000110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1011010000110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1011010000110011010) && ({row_reg, col_reg}<19'b1011010010011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1011010010011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1011010010011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1011010010011101010) && ({row_reg, col_reg}<19'b1011010010011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011010010011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1011010010011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011010010011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1011010010011101111) && ({row_reg, col_reg}<19'b1011010010100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011010010100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1011010010100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1011010010100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1011010010100000100) && ({row_reg, col_reg}<19'b1011010010101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1011010010101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1011010010101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1011010010110000000) && ({row_reg, col_reg}<19'b1011010010110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011010010110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1011010010110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1011010010110011010) && ({row_reg, col_reg}<19'b1011010100011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1011010100011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1011010100011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1011010100011101010) && ({row_reg, col_reg}<19'b1011010100011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011010100011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1011010100011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011010100011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1011010100011101111) && ({row_reg, col_reg}<19'b1011010100100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011010100100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1011010100100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1011010100100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1011010100100000100) && ({row_reg, col_reg}<19'b1011010100101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1011010100101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1011010100101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1011010100110000000) && ({row_reg, col_reg}<19'b1011010100110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011010100110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1011010100110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1011010100110011010) && ({row_reg, col_reg}<19'b1011010110011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1011010110011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1011010110011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1011010110011101010) && ({row_reg, col_reg}<19'b1011010110011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011010110011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1011010110011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011010110011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1011010110011101111) && ({row_reg, col_reg}<19'b1011010110100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011010110100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1011010110100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1011010110100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1011010110100000100) && ({row_reg, col_reg}<19'b1011010110101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1011010110101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1011010110101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1011010110110000000) && ({row_reg, col_reg}<19'b1011010110110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011010110110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1011010110110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1011010110110011010) && ({row_reg, col_reg}<19'b1011011000011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1011011000011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1011011000011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1011011000011101010) && ({row_reg, col_reg}<19'b1011011000011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011011000011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1011011000011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011011000011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1011011000011101111) && ({row_reg, col_reg}<19'b1011011000100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011011000100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1011011000100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1011011000100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1011011000100000100) && ({row_reg, col_reg}<19'b1011011000101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1011011000101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1011011000101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1011011000110000000) && ({row_reg, col_reg}<19'b1011011000110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011011000110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1011011000110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1011011000110011010) && ({row_reg, col_reg}<19'b1011011010011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1011011010011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1011011010011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1011011010011101010) && ({row_reg, col_reg}<19'b1011011010011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011011010011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1011011010011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011011010011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1011011010011101111) && ({row_reg, col_reg}<19'b1011011010100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011011010100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1011011010100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1011011010100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1011011010100000100) && ({row_reg, col_reg}<19'b1011011010101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1011011010101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1011011010101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1011011010110000000) && ({row_reg, col_reg}<19'b1011011010110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011011010110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1011011010110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1011011010110011010) && ({row_reg, col_reg}<19'b1011011100011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1011011100011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1011011100011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1011011100011101010) && ({row_reg, col_reg}<19'b1011011100011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011011100011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1011011100011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011011100011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1011011100011101111) && ({row_reg, col_reg}<19'b1011011100100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011011100100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1011011100100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1011011100100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1011011100100000100) && ({row_reg, col_reg}<19'b1011011100101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1011011100101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1011011100101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1011011100110000000) && ({row_reg, col_reg}<19'b1011011100110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011011100110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1011011100110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1011011100110011010) && ({row_reg, col_reg}<19'b1011011110011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1011011110011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1011011110011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1011011110011101010) && ({row_reg, col_reg}<19'b1011011110011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011011110011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1011011110011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011011110011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1011011110011101111) && ({row_reg, col_reg}<19'b1011011110100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011011110100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1011011110100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1011011110100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1011011110100000100) && ({row_reg, col_reg}<19'b1011011110101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1011011110101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1011011110101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1011011110110000000) && ({row_reg, col_reg}<19'b1011011110110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011011110110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1011011110110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1011011110110011010) && ({row_reg, col_reg}<19'b1011100000011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1011100000011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1011100000011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1011100000011101010) && ({row_reg, col_reg}<19'b1011100000011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011100000011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1011100000011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011100000011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1011100000011101111) && ({row_reg, col_reg}<19'b1011100000100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011100000100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1011100000100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1011100000100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1011100000100000100) && ({row_reg, col_reg}<19'b1011100000101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1011100000101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1011100000101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1011100000110000000) && ({row_reg, col_reg}<19'b1011100000110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011100000110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1011100000110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1011100000110011010) && ({row_reg, col_reg}<19'b1011100010011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1011100010011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1011100010011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1011100010011101010) && ({row_reg, col_reg}<19'b1011100010011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011100010011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1011100010011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011100010011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1011100010011101111) && ({row_reg, col_reg}<19'b1011100010100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011100010100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1011100010100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1011100010100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1011100010100000100) && ({row_reg, col_reg}<19'b1011100010101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1011100010101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1011100010101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1011100010110000000) && ({row_reg, col_reg}<19'b1011100010110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011100010110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1011100010110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1011100010110011010) && ({row_reg, col_reg}<19'b1011100100011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1011100100011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1011100100011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1011100100011101010) && ({row_reg, col_reg}<19'b1011100100011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011100100011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1011100100011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011100100011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1011100100011101111) && ({row_reg, col_reg}<19'b1011100100100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011100100100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1011100100100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1011100100100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1011100100100000100) && ({row_reg, col_reg}<19'b1011100100101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1011100100101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1011100100101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1011100100110000000) && ({row_reg, col_reg}<19'b1011100100110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011100100110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1011100100110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1011100100110011010) && ({row_reg, col_reg}<19'b1011100110011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1011100110011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1011100110011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1011100110011101010) && ({row_reg, col_reg}<19'b1011100110011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011100110011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1011100110011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011100110011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1011100110011101111) && ({row_reg, col_reg}<19'b1011100110100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011100110100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1011100110100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1011100110100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1011100110100000100) && ({row_reg, col_reg}<19'b1011100110101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1011100110101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1011100110101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1011100110110000000) && ({row_reg, col_reg}<19'b1011100110110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011100110110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1011100110110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1011100110110011010) && ({row_reg, col_reg}<19'b1011101000011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1011101000011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1011101000011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1011101000011101010) && ({row_reg, col_reg}<19'b1011101000011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011101000011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1011101000011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011101000011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1011101000011101111) && ({row_reg, col_reg}<19'b1011101000100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011101000100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1011101000100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1011101000100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1011101000100000100) && ({row_reg, col_reg}<19'b1011101000101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1011101000101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1011101000101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1011101000110000000) && ({row_reg, col_reg}<19'b1011101000110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011101000110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1011101000110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1011101000110011010) && ({row_reg, col_reg}<19'b1011101010011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1011101010011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1011101010011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1011101010011101010) && ({row_reg, col_reg}<19'b1011101010011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011101010011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1011101010011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011101010011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1011101010011101111) && ({row_reg, col_reg}<19'b1011101010100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011101010100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1011101010100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1011101010100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1011101010100000100) && ({row_reg, col_reg}<19'b1011101010101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1011101010101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1011101010101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1011101010110000000) && ({row_reg, col_reg}<19'b1011101010110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011101010110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1011101010110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1011101010110011010) && ({row_reg, col_reg}<19'b1011101100011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1011101100011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1011101100011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1011101100011101010) && ({row_reg, col_reg}<19'b1011101100011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011101100011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1011101100011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011101100011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1011101100011101111) && ({row_reg, col_reg}<19'b1011101100100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011101100100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1011101100100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1011101100100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1011101100100000100) && ({row_reg, col_reg}<19'b1011101100101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1011101100101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1011101100101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1011101100110000000) && ({row_reg, col_reg}<19'b1011101100110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011101100110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1011101100110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1011101100110011010) && ({row_reg, col_reg}<19'b1011101110011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1011101110011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1011101110011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1011101110011101010) && ({row_reg, col_reg}<19'b1011101110011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011101110011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1011101110011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011101110011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1011101110011101111) && ({row_reg, col_reg}<19'b1011101110100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011101110100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1011101110100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1011101110100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1011101110100000100) && ({row_reg, col_reg}<19'b1011101110101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1011101110101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1011101110101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1011101110110000000) && ({row_reg, col_reg}<19'b1011101110110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011101110110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1011101110110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1011101110110011010) && ({row_reg, col_reg}<19'b1011110000011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1011110000011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1011110000011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1011110000011101010) && ({row_reg, col_reg}<19'b1011110000011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011110000011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1011110000011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011110000011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1011110000011101111) && ({row_reg, col_reg}<19'b1011110000100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011110000100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1011110000100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1011110000100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1011110000100000100) && ({row_reg, col_reg}<19'b1011110000101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1011110000101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1011110000101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1011110000110000000) && ({row_reg, col_reg}<19'b1011110000110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011110000110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1011110000110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1011110000110011010) && ({row_reg, col_reg}<19'b1011110010011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1011110010011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1011110010011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1011110010011101010) && ({row_reg, col_reg}<19'b1011110010011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011110010011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1011110010011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011110010011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1011110010011101111) && ({row_reg, col_reg}<19'b1011110010100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011110010100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1011110010100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1011110010100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1011110010100000100) && ({row_reg, col_reg}<19'b1011110010101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1011110010101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1011110010101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1011110010110000000) && ({row_reg, col_reg}<19'b1011110010110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011110010110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1011110010110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1011110010110011010) && ({row_reg, col_reg}<19'b1011110100011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1011110100011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1011110100011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1011110100011101010) && ({row_reg, col_reg}<19'b1011110100011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011110100011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1011110100011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011110100011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1011110100011101111) && ({row_reg, col_reg}<19'b1011110100100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011110100100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1011110100100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1011110100100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1011110100100000100) && ({row_reg, col_reg}<19'b1011110100101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1011110100101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1011110100101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1011110100110000000) && ({row_reg, col_reg}<19'b1011110100110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011110100110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1011110100110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1011110100110011010) && ({row_reg, col_reg}<19'b1011110110011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1011110110011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1011110110011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1011110110011101010) && ({row_reg, col_reg}<19'b1011110110011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011110110011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1011110110011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011110110011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1011110110011101111) && ({row_reg, col_reg}<19'b1011110110100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011110110100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1011110110100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1011110110100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1011110110100000100) && ({row_reg, col_reg}<19'b1011110110101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1011110110101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1011110110101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1011110110110000000) && ({row_reg, col_reg}<19'b1011110110110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011110110110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1011110110110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1011110110110011010) && ({row_reg, col_reg}<19'b1011111000011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1011111000011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1011111000011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1011111000011101010) && ({row_reg, col_reg}<19'b1011111000011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011111000011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1011111000011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011111000011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1011111000011101111) && ({row_reg, col_reg}<19'b1011111000100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011111000100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1011111000100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1011111000100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1011111000100000100) && ({row_reg, col_reg}<19'b1011111000101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1011111000101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1011111000101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1011111000110000000) && ({row_reg, col_reg}<19'b1011111000110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011111000110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1011111000110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1011111000110011010) && ({row_reg, col_reg}<19'b1011111010011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1011111010011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1011111010011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1011111010011101010) && ({row_reg, col_reg}<19'b1011111010011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011111010011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1011111010011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011111010011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1011111010011101111) && ({row_reg, col_reg}<19'b1011111010100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011111010100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1011111010100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1011111010100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1011111010100000100) && ({row_reg, col_reg}<19'b1011111010101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1011111010101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1011111010101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1011111010110000000) && ({row_reg, col_reg}<19'b1011111010110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011111010110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1011111010110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1011111010110011010) && ({row_reg, col_reg}<19'b1011111100011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1011111100011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1011111100011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1011111100011101010) && ({row_reg, col_reg}<19'b1011111100011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011111100011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1011111100011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011111100011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1011111100011101111) && ({row_reg, col_reg}<19'b1011111100100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011111100100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1011111100100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1011111100100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1011111100100000100) && ({row_reg, col_reg}<19'b1011111100101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1011111100101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1011111100101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1011111100110000000) && ({row_reg, col_reg}<19'b1011111100110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011111100110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1011111100110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1011111100110011010) && ({row_reg, col_reg}<19'b1011111110011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1011111110011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1011111110011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1011111110011101010) && ({row_reg, col_reg}<19'b1011111110011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011111110011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1011111110011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011111110011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1011111110011101111) && ({row_reg, col_reg}<19'b1011111110100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011111110100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1011111110100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1011111110100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1011111110100000100) && ({row_reg, col_reg}<19'b1011111110101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1011111110101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1011111110101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1011111110110000000) && ({row_reg, col_reg}<19'b1011111110110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011111110110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1011111110110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1011111110110011010) && ({row_reg, col_reg}<19'b1100000000011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1100000000011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1100000000011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1100000000011101010) && ({row_reg, col_reg}<19'b1100000000011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100000000011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1100000000011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100000000011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1100000000011101111) && ({row_reg, col_reg}<19'b1100000000100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100000000100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1100000000100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1100000000100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1100000000100000100) && ({row_reg, col_reg}<19'b1100000000101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1100000000101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1100000000101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1100000000110000000) && ({row_reg, col_reg}<19'b1100000000110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100000000110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1100000000110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1100000000110011010) && ({row_reg, col_reg}<19'b1100000010011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1100000010011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1100000010011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1100000010011101010) && ({row_reg, col_reg}<19'b1100000010011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100000010011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1100000010011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100000010011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1100000010011101111) && ({row_reg, col_reg}<19'b1100000010100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100000010100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1100000010100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1100000010100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1100000010100000100) && ({row_reg, col_reg}<19'b1100000010101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1100000010101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1100000010101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1100000010110000000) && ({row_reg, col_reg}<19'b1100000010110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100000010110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1100000010110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1100000010110011010) && ({row_reg, col_reg}<19'b1100000100011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1100000100011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1100000100011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1100000100011101010) && ({row_reg, col_reg}<19'b1100000100011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100000100011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1100000100011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100000100011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1100000100011101111) && ({row_reg, col_reg}<19'b1100000100100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100000100100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1100000100100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1100000100100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1100000100100000100) && ({row_reg, col_reg}<19'b1100000100101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1100000100101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1100000100101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1100000100110000000) && ({row_reg, col_reg}<19'b1100000100110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100000100110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1100000100110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1100000100110011010) && ({row_reg, col_reg}<19'b1100000110011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1100000110011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1100000110011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1100000110011101010) && ({row_reg, col_reg}<19'b1100000110011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100000110011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1100000110011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100000110011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1100000110011101111) && ({row_reg, col_reg}<19'b1100000110100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100000110100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1100000110100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1100000110100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1100000110100000100) && ({row_reg, col_reg}<19'b1100000110101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1100000110101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1100000110101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1100000110110000000) && ({row_reg, col_reg}<19'b1100000110110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100000110110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1100000110110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1100000110110011010) && ({row_reg, col_reg}<19'b1100001000011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1100001000011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1100001000011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1100001000011101010) && ({row_reg, col_reg}<19'b1100001000011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100001000011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1100001000011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100001000011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1100001000011101111) && ({row_reg, col_reg}<19'b1100001000100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100001000100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1100001000100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1100001000100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1100001000100000100) && ({row_reg, col_reg}<19'b1100001000101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1100001000101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1100001000101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1100001000110000000) && ({row_reg, col_reg}<19'b1100001000110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100001000110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1100001000110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1100001000110011010) && ({row_reg, col_reg}<19'b1100001010011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1100001010011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1100001010011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1100001010011101010) && ({row_reg, col_reg}<19'b1100001010011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100001010011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1100001010011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100001010011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1100001010011101111) && ({row_reg, col_reg}<19'b1100001010100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100001010100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1100001010100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1100001010100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1100001010100000100) && ({row_reg, col_reg}<19'b1100001010101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1100001010101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1100001010101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1100001010110000000) && ({row_reg, col_reg}<19'b1100001010110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100001010110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1100001010110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1100001010110011010) && ({row_reg, col_reg}<19'b1100001100011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1100001100011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1100001100011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1100001100011101010) && ({row_reg, col_reg}<19'b1100001100011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100001100011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1100001100011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100001100011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1100001100011101111) && ({row_reg, col_reg}<19'b1100001100100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100001100100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1100001100100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1100001100100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1100001100100000100) && ({row_reg, col_reg}<19'b1100001100101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1100001100101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1100001100101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1100001100110000000) && ({row_reg, col_reg}<19'b1100001100110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100001100110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1100001100110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1100001100110011010) && ({row_reg, col_reg}<19'b1100001110011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1100001110011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1100001110011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1100001110011101010) && ({row_reg, col_reg}<19'b1100001110011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100001110011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1100001110011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100001110011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1100001110011101111) && ({row_reg, col_reg}<19'b1100001110100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100001110100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1100001110100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1100001110100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1100001110100000100) && ({row_reg, col_reg}<19'b1100001110101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1100001110101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1100001110101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1100001110110000000) && ({row_reg, col_reg}<19'b1100001110110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100001110110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1100001110110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1100001110110011010) && ({row_reg, col_reg}<19'b1100010000011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1100010000011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1100010000011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1100010000011101010) && ({row_reg, col_reg}<19'b1100010000011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100010000011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1100010000011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100010000011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1100010000011101111) && ({row_reg, col_reg}<19'b1100010000100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100010000100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1100010000100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1100010000100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1100010000100000100) && ({row_reg, col_reg}<19'b1100010000101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1100010000101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1100010000101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1100010000110000000) && ({row_reg, col_reg}<19'b1100010000110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100010000110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1100010000110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1100010000110011010) && ({row_reg, col_reg}<19'b1100010010011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1100010010011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1100010010011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1100010010011101010) && ({row_reg, col_reg}<19'b1100010010011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100010010011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1100010010011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100010010011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1100010010011101111) && ({row_reg, col_reg}<19'b1100010010100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100010010100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1100010010100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1100010010100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1100010010100000100) && ({row_reg, col_reg}<19'b1100010010101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1100010010101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1100010010101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1100010010110000000) && ({row_reg, col_reg}<19'b1100010010110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100010010110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1100010010110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1100010010110011010) && ({row_reg, col_reg}<19'b1100010100011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1100010100011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1100010100011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1100010100011101010) && ({row_reg, col_reg}<19'b1100010100011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100010100011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1100010100011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100010100011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1100010100011101111) && ({row_reg, col_reg}<19'b1100010100100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100010100100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1100010100100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1100010100100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1100010100100000100) && ({row_reg, col_reg}<19'b1100010100101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1100010100101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1100010100101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1100010100110000000) && ({row_reg, col_reg}<19'b1100010100110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100010100110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1100010100110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1100010100110011010) && ({row_reg, col_reg}<19'b1100010110011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1100010110011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1100010110011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1100010110011101010) && ({row_reg, col_reg}<19'b1100010110011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100010110011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1100010110011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100010110011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1100010110011101111) && ({row_reg, col_reg}<19'b1100010110100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100010110100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1100010110100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1100010110100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1100010110100000100) && ({row_reg, col_reg}<19'b1100010110101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1100010110101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1100010110101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1100010110110000000) && ({row_reg, col_reg}<19'b1100010110110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100010110110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1100010110110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1100010110110011010) && ({row_reg, col_reg}<19'b1100011000011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1100011000011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1100011000011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1100011000011101010) && ({row_reg, col_reg}<19'b1100011000011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100011000011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1100011000011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100011000011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1100011000011101111) && ({row_reg, col_reg}<19'b1100011000100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100011000100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1100011000100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1100011000100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1100011000100000100) && ({row_reg, col_reg}<19'b1100011000101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1100011000101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1100011000101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1100011000110000000) && ({row_reg, col_reg}<19'b1100011000110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100011000110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1100011000110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1100011000110011010) && ({row_reg, col_reg}<19'b1100011010011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1100011010011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1100011010011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1100011010011101010) && ({row_reg, col_reg}<19'b1100011010011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100011010011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1100011010011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100011010011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1100011010011101111) && ({row_reg, col_reg}<19'b1100011010100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100011010100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1100011010100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1100011010100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1100011010100000100) && ({row_reg, col_reg}<19'b1100011010101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1100011010101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1100011010101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1100011010110000000) && ({row_reg, col_reg}<19'b1100011010110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100011010110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1100011010110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1100011010110011010) && ({row_reg, col_reg}<19'b1100011100011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1100011100011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1100011100011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1100011100011101010) && ({row_reg, col_reg}<19'b1100011100011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100011100011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1100011100011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100011100011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1100011100011101111) && ({row_reg, col_reg}<19'b1100011100100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100011100100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1100011100100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1100011100100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1100011100100000100) && ({row_reg, col_reg}<19'b1100011100101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1100011100101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1100011100101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1100011100110000000) && ({row_reg, col_reg}<19'b1100011100110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100011100110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1100011100110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1100011100110011010) && ({row_reg, col_reg}<19'b1100011110011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1100011110011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1100011110011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1100011110011101010) && ({row_reg, col_reg}<19'b1100011110011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100011110011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1100011110011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100011110011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1100011110011101111) && ({row_reg, col_reg}<19'b1100011110100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100011110100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1100011110100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1100011110100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1100011110100000100) && ({row_reg, col_reg}<19'b1100011110101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1100011110101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1100011110101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1100011110110000000) && ({row_reg, col_reg}<19'b1100011110110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100011110110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1100011110110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1100011110110011010) && ({row_reg, col_reg}<19'b1100100000011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1100100000011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1100100000011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1100100000011101010) && ({row_reg, col_reg}<19'b1100100000011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100100000011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1100100000011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100100000011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1100100000011101111) && ({row_reg, col_reg}<19'b1100100000100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100100000100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1100100000100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1100100000100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1100100000100000100) && ({row_reg, col_reg}<19'b1100100000101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1100100000101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1100100000101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1100100000110000000) && ({row_reg, col_reg}<19'b1100100000110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100100000110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1100100000110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1100100000110011010) && ({row_reg, col_reg}<19'b1100100010011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1100100010011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1100100010011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1100100010011101010) && ({row_reg, col_reg}<19'b1100100010011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100100010011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1100100010011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100100010011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1100100010011101111) && ({row_reg, col_reg}<19'b1100100010100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100100010100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1100100010100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1100100010100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1100100010100000100) && ({row_reg, col_reg}<19'b1100100010101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1100100010101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1100100010101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1100100010110000000) && ({row_reg, col_reg}<19'b1100100010110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100100010110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1100100010110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1100100010110011010) && ({row_reg, col_reg}<19'b1100100100011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1100100100011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1100100100011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1100100100011101010) && ({row_reg, col_reg}<19'b1100100100011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100100100011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1100100100011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100100100011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1100100100011101111) && ({row_reg, col_reg}<19'b1100100100100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100100100100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1100100100100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1100100100100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1100100100100000100) && ({row_reg, col_reg}<19'b1100100100101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1100100100101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1100100100101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1100100100110000000) && ({row_reg, col_reg}<19'b1100100100110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100100100110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1100100100110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1100100100110011010) && ({row_reg, col_reg}<19'b1100100110011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1100100110011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1100100110011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1100100110011101010) && ({row_reg, col_reg}<19'b1100100110011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100100110011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1100100110011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100100110011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1100100110011101111) && ({row_reg, col_reg}<19'b1100100110100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100100110100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1100100110100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1100100110100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1100100110100000100) && ({row_reg, col_reg}<19'b1100100110101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1100100110101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1100100110101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1100100110110000000) && ({row_reg, col_reg}<19'b1100100110110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100100110110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1100100110110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1100100110110011010) && ({row_reg, col_reg}<19'b1100101000011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1100101000011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1100101000011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1100101000011101010) && ({row_reg, col_reg}<19'b1100101000011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100101000011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1100101000011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100101000011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1100101000011101111) && ({row_reg, col_reg}<19'b1100101000100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100101000100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1100101000100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1100101000100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1100101000100000100) && ({row_reg, col_reg}<19'b1100101000101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1100101000101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1100101000101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1100101000110000000) && ({row_reg, col_reg}<19'b1100101000110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100101000110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1100101000110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1100101000110011010) && ({row_reg, col_reg}<19'b1100101010011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1100101010011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1100101010011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1100101010011101010) && ({row_reg, col_reg}<19'b1100101010011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100101010011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1100101010011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100101010011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1100101010011101111) && ({row_reg, col_reg}<19'b1100101010100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100101010100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1100101010100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1100101010100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1100101010100000100) && ({row_reg, col_reg}<19'b1100101010101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1100101010101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1100101010101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1100101010110000000) && ({row_reg, col_reg}<19'b1100101010110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100101010110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1100101010110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1100101010110011010) && ({row_reg, col_reg}<19'b1100101100011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1100101100011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1100101100011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1100101100011101010) && ({row_reg, col_reg}<19'b1100101100011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100101100011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1100101100011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100101100011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1100101100011101111) && ({row_reg, col_reg}<19'b1100101100100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100101100100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1100101100100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1100101100100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1100101100100000100) && ({row_reg, col_reg}<19'b1100101100101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1100101100101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1100101100101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1100101100110000000) && ({row_reg, col_reg}<19'b1100101100110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100101100110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1100101100110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1100101100110011010) && ({row_reg, col_reg}<19'b1100101110011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1100101110011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1100101110011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1100101110011101010) && ({row_reg, col_reg}<19'b1100101110011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100101110011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1100101110011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100101110011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1100101110011101111) && ({row_reg, col_reg}<19'b1100101110100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100101110100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1100101110100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1100101110100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1100101110100000100) && ({row_reg, col_reg}<19'b1100101110101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1100101110101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1100101110101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1100101110110000000) && ({row_reg, col_reg}<19'b1100101110110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100101110110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1100101110110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1100101110110011010) && ({row_reg, col_reg}<19'b1100110000011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1100110000011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1100110000011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1100110000011101010) && ({row_reg, col_reg}<19'b1100110000011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100110000011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1100110000011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100110000011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1100110000011101111) && ({row_reg, col_reg}<19'b1100110000100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100110000100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1100110000100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1100110000100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1100110000100000100) && ({row_reg, col_reg}<19'b1100110000101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1100110000101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1100110000101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1100110000110000000) && ({row_reg, col_reg}<19'b1100110000110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100110000110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1100110000110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1100110000110011010) && ({row_reg, col_reg}<19'b1100110010011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1100110010011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1100110010011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1100110010011101010) && ({row_reg, col_reg}<19'b1100110010011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100110010011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1100110010011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100110010011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1100110010011101111) && ({row_reg, col_reg}<19'b1100110010100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100110010100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1100110010100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1100110010100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1100110010100000100) && ({row_reg, col_reg}<19'b1100110010101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1100110010101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1100110010101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1100110010110000000) && ({row_reg, col_reg}<19'b1100110010110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100110010110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1100110010110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1100110010110011010) && ({row_reg, col_reg}<19'b1100110100011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1100110100011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1100110100011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1100110100011101010) && ({row_reg, col_reg}<19'b1100110100011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100110100011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1100110100011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100110100011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1100110100011101111) && ({row_reg, col_reg}<19'b1100110100100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100110100100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1100110100100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1100110100100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1100110100100000100) && ({row_reg, col_reg}<19'b1100110100101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1100110100101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1100110100101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1100110100110000000) && ({row_reg, col_reg}<19'b1100110100110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100110100110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1100110100110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1100110100110011010) && ({row_reg, col_reg}<19'b1100110110011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1100110110011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1100110110011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1100110110011101010) && ({row_reg, col_reg}<19'b1100110110011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100110110011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1100110110011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100110110011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1100110110011101111) && ({row_reg, col_reg}<19'b1100110110100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100110110100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1100110110100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1100110110100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1100110110100000100) && ({row_reg, col_reg}<19'b1100110110101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1100110110101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1100110110101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1100110110110000000) && ({row_reg, col_reg}<19'b1100110110110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100110110110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1100110110110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1100110110110011010) && ({row_reg, col_reg}<19'b1100111000011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1100111000011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1100111000011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1100111000011101010) && ({row_reg, col_reg}<19'b1100111000011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100111000011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1100111000011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100111000011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1100111000011101111) && ({row_reg, col_reg}<19'b1100111000100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100111000100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1100111000100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1100111000100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1100111000100000100) && ({row_reg, col_reg}<19'b1100111000101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1100111000101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1100111000101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1100111000110000000) && ({row_reg, col_reg}<19'b1100111000110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100111000110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1100111000110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1100111000110011010) && ({row_reg, col_reg}<19'b1100111010011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1100111010011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1100111010011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1100111010011101010) && ({row_reg, col_reg}<19'b1100111010011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100111010011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1100111010011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100111010011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1100111010011101111) && ({row_reg, col_reg}<19'b1100111010100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100111010100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1100111010100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1100111010100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1100111010100000100) && ({row_reg, col_reg}<19'b1100111010101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1100111010101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1100111010101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1100111010110000000) && ({row_reg, col_reg}<19'b1100111010110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100111010110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1100111010110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1100111010110011010) && ({row_reg, col_reg}<19'b1100111100011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1100111100011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1100111100011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1100111100011101010) && ({row_reg, col_reg}<19'b1100111100011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100111100011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1100111100011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100111100011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1100111100011101111) && ({row_reg, col_reg}<19'b1100111100100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100111100100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1100111100100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1100111100100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1100111100100000100) && ({row_reg, col_reg}<19'b1100111100101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1100111100101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1100111100101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1100111100110000000) && ({row_reg, col_reg}<19'b1100111100110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100111100110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1100111100110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1100111100110011010) && ({row_reg, col_reg}<19'b1100111110011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1100111110011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1100111110011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1100111110011101010) && ({row_reg, col_reg}<19'b1100111110011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100111110011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1100111110011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100111110011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1100111110011101111) && ({row_reg, col_reg}<19'b1100111110100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100111110100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1100111110100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1100111110100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1100111110100000100) && ({row_reg, col_reg}<19'b1100111110101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1100111110101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1100111110101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1100111110110000000) && ({row_reg, col_reg}<19'b1100111110110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100111110110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1100111110110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1100111110110011010) && ({row_reg, col_reg}<19'b1101000000011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1101000000011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1101000000011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1101000000011101010) && ({row_reg, col_reg}<19'b1101000000011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101000000011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1101000000011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101000000011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1101000000011101111) && ({row_reg, col_reg}<19'b1101000000100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101000000100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1101000000100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1101000000100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1101000000100000100) && ({row_reg, col_reg}<19'b1101000000101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1101000000101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1101000000101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1101000000110000000) && ({row_reg, col_reg}<19'b1101000000110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101000000110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1101000000110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1101000000110011010) && ({row_reg, col_reg}<19'b1101000010011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1101000010011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1101000010011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1101000010011101010) && ({row_reg, col_reg}<19'b1101000010011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101000010011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1101000010011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101000010011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1101000010011101111) && ({row_reg, col_reg}<19'b1101000010100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101000010100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1101000010100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1101000010100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1101000010100000100) && ({row_reg, col_reg}<19'b1101000010101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1101000010101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1101000010101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1101000010110000000) && ({row_reg, col_reg}<19'b1101000010110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101000010110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1101000010110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1101000010110011010) && ({row_reg, col_reg}<19'b1101000100011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1101000100011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1101000100011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1101000100011101010) && ({row_reg, col_reg}<19'b1101000100011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101000100011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1101000100011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101000100011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1101000100011101111) && ({row_reg, col_reg}<19'b1101000100100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101000100100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1101000100100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1101000100100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1101000100100000100) && ({row_reg, col_reg}<19'b1101000100101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1101000100101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1101000100101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1101000100110000000) && ({row_reg, col_reg}<19'b1101000100110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101000100110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1101000100110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1101000100110011010) && ({row_reg, col_reg}<19'b1101000110011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1101000110011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1101000110011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1101000110011101010) && ({row_reg, col_reg}<19'b1101000110011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101000110011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1101000110011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101000110011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1101000110011101111) && ({row_reg, col_reg}<19'b1101000110100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101000110100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1101000110100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1101000110100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1101000110100000100) && ({row_reg, col_reg}<19'b1101000110101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1101000110101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1101000110101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1101000110110000000) && ({row_reg, col_reg}<19'b1101000110110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101000110110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1101000110110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1101000110110011010) && ({row_reg, col_reg}<19'b1101001000011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1101001000011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1101001000011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1101001000011101010) && ({row_reg, col_reg}<19'b1101001000011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101001000011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1101001000011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101001000011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1101001000011101111) && ({row_reg, col_reg}<19'b1101001000100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101001000100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1101001000100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1101001000100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1101001000100000100) && ({row_reg, col_reg}<19'b1101001000101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1101001000101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1101001000101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1101001000110000000) && ({row_reg, col_reg}<19'b1101001000110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101001000110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1101001000110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1101001000110011010) && ({row_reg, col_reg}<19'b1101001010011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1101001010011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1101001010011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1101001010011101010) && ({row_reg, col_reg}<19'b1101001010011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101001010011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1101001010011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101001010011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1101001010011101111) && ({row_reg, col_reg}<19'b1101001010100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101001010100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1101001010100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1101001010100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1101001010100000100) && ({row_reg, col_reg}<19'b1101001010101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1101001010101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1101001010101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1101001010110000000) && ({row_reg, col_reg}<19'b1101001010110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101001010110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1101001010110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1101001010110011010) && ({row_reg, col_reg}<19'b1101001100011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1101001100011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1101001100011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1101001100011101010) && ({row_reg, col_reg}<19'b1101001100011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101001100011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1101001100011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101001100011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1101001100011101111) && ({row_reg, col_reg}<19'b1101001100100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101001100100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1101001100100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1101001100100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1101001100100000100) && ({row_reg, col_reg}<19'b1101001100101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1101001100101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1101001100101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1101001100110000000) && ({row_reg, col_reg}<19'b1101001100110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101001100110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1101001100110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1101001100110011010) && ({row_reg, col_reg}<19'b1101001110011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1101001110011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1101001110011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1101001110011101010) && ({row_reg, col_reg}<19'b1101001110011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101001110011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1101001110011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101001110011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1101001110011101111) && ({row_reg, col_reg}<19'b1101001110100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101001110100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1101001110100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1101001110100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1101001110100000100) && ({row_reg, col_reg}<19'b1101001110101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1101001110101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1101001110101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1101001110110000000) && ({row_reg, col_reg}<19'b1101001110110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101001110110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1101001110110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1101001110110011010) && ({row_reg, col_reg}<19'b1101010000011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1101010000011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1101010000011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1101010000011101010) && ({row_reg, col_reg}<19'b1101010000011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101010000011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1101010000011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101010000011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1101010000011101111) && ({row_reg, col_reg}<19'b1101010000100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101010000100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1101010000100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1101010000100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1101010000100000100) && ({row_reg, col_reg}<19'b1101010000101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1101010000101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1101010000101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1101010000110000000) && ({row_reg, col_reg}<19'b1101010000110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101010000110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1101010000110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1101010000110011010) && ({row_reg, col_reg}<19'b1101010010011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1101010010011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1101010010011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1101010010011101010) && ({row_reg, col_reg}<19'b1101010010011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101010010011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1101010010011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101010010011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1101010010011101111) && ({row_reg, col_reg}<19'b1101010010100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101010010100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1101010010100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1101010010100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1101010010100000100) && ({row_reg, col_reg}<19'b1101010010101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1101010010101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1101010010101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1101010010110000000) && ({row_reg, col_reg}<19'b1101010010110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101010010110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1101010010110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1101010010110011010) && ({row_reg, col_reg}<19'b1101010100011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1101010100011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1101010100011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1101010100011101010) && ({row_reg, col_reg}<19'b1101010100011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101010100011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1101010100011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101010100011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1101010100011101111) && ({row_reg, col_reg}<19'b1101010100100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101010100100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1101010100100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1101010100100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1101010100100000100) && ({row_reg, col_reg}<19'b1101010100101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1101010100101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1101010100101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1101010100110000000) && ({row_reg, col_reg}<19'b1101010100110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101010100110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1101010100110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1101010100110011010) && ({row_reg, col_reg}<19'b1101010110011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1101010110011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1101010110011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1101010110011101010) && ({row_reg, col_reg}<19'b1101010110011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101010110011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1101010110011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101010110011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1101010110011101111) && ({row_reg, col_reg}<19'b1101010110100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101010110100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1101010110100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1101010110100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1101010110100000100) && ({row_reg, col_reg}<19'b1101010110101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1101010110101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1101010110101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1101010110110000000) && ({row_reg, col_reg}<19'b1101010110110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101010110110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1101010110110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1101010110110011010) && ({row_reg, col_reg}<19'b1101011000011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1101011000011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1101011000011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1101011000011101010) && ({row_reg, col_reg}<19'b1101011000011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101011000011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1101011000011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101011000011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1101011000011101111) && ({row_reg, col_reg}<19'b1101011000100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101011000100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1101011000100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1101011000100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1101011000100000100) && ({row_reg, col_reg}<19'b1101011000101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1101011000101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1101011000101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1101011000110000000) && ({row_reg, col_reg}<19'b1101011000110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101011000110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1101011000110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1101011000110011010) && ({row_reg, col_reg}<19'b1101011010011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1101011010011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1101011010011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1101011010011101010) && ({row_reg, col_reg}<19'b1101011010011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101011010011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1101011010011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101011010011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1101011010011101111) && ({row_reg, col_reg}<19'b1101011010100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101011010100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1101011010100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1101011010100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1101011010100000100) && ({row_reg, col_reg}<19'b1101011010101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1101011010101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1101011010101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1101011010110000000) && ({row_reg, col_reg}<19'b1101011010110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101011010110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1101011010110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1101011010110011010) && ({row_reg, col_reg}<19'b1101011100011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1101011100011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1101011100011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1101011100011101010) && ({row_reg, col_reg}<19'b1101011100011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101011100011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1101011100011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101011100011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1101011100011101111) && ({row_reg, col_reg}<19'b1101011100100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101011100100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1101011100100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1101011100100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1101011100100000100) && ({row_reg, col_reg}<19'b1101011100101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1101011100101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1101011100101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1101011100110000000) && ({row_reg, col_reg}<19'b1101011100110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101011100110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1101011100110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1101011100110011010) && ({row_reg, col_reg}<19'b1101011110011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1101011110011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1101011110011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1101011110011101010) && ({row_reg, col_reg}<19'b1101011110011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101011110011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1101011110011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101011110011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1101011110011101111) && ({row_reg, col_reg}<19'b1101011110100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101011110100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1101011110100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1101011110100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1101011110100000100) && ({row_reg, col_reg}<19'b1101011110101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1101011110101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1101011110101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1101011110110000000) && ({row_reg, col_reg}<19'b1101011110110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101011110110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1101011110110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1101011110110011010) && ({row_reg, col_reg}<19'b1101100000011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1101100000011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1101100000011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1101100000011101010) && ({row_reg, col_reg}<19'b1101100000011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101100000011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1101100000011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101100000011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1101100000011101111) && ({row_reg, col_reg}<19'b1101100000100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101100000100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1101100000100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1101100000100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1101100000100000100) && ({row_reg, col_reg}<19'b1101100000101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1101100000101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1101100000101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1101100000110000000) && ({row_reg, col_reg}<19'b1101100000110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101100000110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1101100000110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1101100000110011010) && ({row_reg, col_reg}<19'b1101100010011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1101100010011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1101100010011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1101100010011101010) && ({row_reg, col_reg}<19'b1101100010011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101100010011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1101100010011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101100010011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1101100010011101111) && ({row_reg, col_reg}<19'b1101100010100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101100010100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1101100010100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1101100010100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1101100010100000100) && ({row_reg, col_reg}<19'b1101100010101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1101100010101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1101100010101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1101100010110000000) && ({row_reg, col_reg}<19'b1101100010110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101100010110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1101100010110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1101100010110011010) && ({row_reg, col_reg}<19'b1101100100011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1101100100011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1101100100011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1101100100011101010) && ({row_reg, col_reg}<19'b1101100100011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101100100011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1101100100011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101100100011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1101100100011101111) && ({row_reg, col_reg}<19'b1101100100100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101100100100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1101100100100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1101100100100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1101100100100000100) && ({row_reg, col_reg}<19'b1101100100101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1101100100101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1101100100101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1101100100110000000) && ({row_reg, col_reg}<19'b1101100100110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101100100110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1101100100110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1101100100110011010) && ({row_reg, col_reg}<19'b1101100110011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1101100110011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1101100110011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1101100110011101010) && ({row_reg, col_reg}<19'b1101100110011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101100110011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1101100110011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101100110011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1101100110011101111) && ({row_reg, col_reg}<19'b1101100110100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101100110100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1101100110100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1101100110100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1101100110100000100) && ({row_reg, col_reg}<19'b1101100110101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1101100110101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1101100110101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1101100110110000000) && ({row_reg, col_reg}<19'b1101100110110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101100110110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1101100110110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1101100110110011010) && ({row_reg, col_reg}<19'b1101101000011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1101101000011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1101101000011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1101101000011101010) && ({row_reg, col_reg}<19'b1101101000011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101101000011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1101101000011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101101000011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1101101000011101111) && ({row_reg, col_reg}<19'b1101101000100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101101000100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1101101000100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1101101000100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1101101000100000100) && ({row_reg, col_reg}<19'b1101101000101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1101101000101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1101101000101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1101101000110000000) && ({row_reg, col_reg}<19'b1101101000110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101101000110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1101101000110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1101101000110011010) && ({row_reg, col_reg}<19'b1101101010011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1101101010011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1101101010011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1101101010011101010) && ({row_reg, col_reg}<19'b1101101010011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101101010011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1101101010011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101101010011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1101101010011101111) && ({row_reg, col_reg}<19'b1101101010100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101101010100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1101101010100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1101101010100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1101101010100000100) && ({row_reg, col_reg}<19'b1101101010101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1101101010101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1101101010101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1101101010110000000) && ({row_reg, col_reg}<19'b1101101010110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101101010110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1101101010110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1101101010110011010) && ({row_reg, col_reg}<19'b1101101100011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1101101100011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1101101100011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1101101100011101010) && ({row_reg, col_reg}<19'b1101101100011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101101100011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1101101100011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101101100011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1101101100011101111) && ({row_reg, col_reg}<19'b1101101100100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101101100100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1101101100100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1101101100100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1101101100100000100) && ({row_reg, col_reg}<19'b1101101100101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1101101100101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1101101100101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1101101100110000000) && ({row_reg, col_reg}<19'b1101101100110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101101100110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1101101100110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1101101100110011010) && ({row_reg, col_reg}<19'b1101101110011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1101101110011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1101101110011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1101101110011101010) && ({row_reg, col_reg}<19'b1101101110011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101101110011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1101101110011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101101110011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1101101110011101111) && ({row_reg, col_reg}<19'b1101101110100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101101110100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1101101110100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1101101110100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1101101110100000100) && ({row_reg, col_reg}<19'b1101101110101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1101101110101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1101101110101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1101101110110000000) && ({row_reg, col_reg}<19'b1101101110110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101101110110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1101101110110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1101101110110011010) && ({row_reg, col_reg}<19'b1101110000011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1101110000011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1101110000011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1101110000011101010) && ({row_reg, col_reg}<19'b1101110000011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101110000011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1101110000011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101110000011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1101110000011101111) && ({row_reg, col_reg}<19'b1101110000100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101110000100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1101110000100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1101110000100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1101110000100000100) && ({row_reg, col_reg}<19'b1101110000101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1101110000101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1101110000101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1101110000110000000) && ({row_reg, col_reg}<19'b1101110000110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101110000110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1101110000110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1101110000110011010) && ({row_reg, col_reg}<19'b1101110010011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1101110010011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1101110010011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1101110010011101010) && ({row_reg, col_reg}<19'b1101110010011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101110010011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1101110010011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101110010011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1101110010011101111) && ({row_reg, col_reg}<19'b1101110010100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101110010100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1101110010100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1101110010100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1101110010100000100) && ({row_reg, col_reg}<19'b1101110010101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1101110010101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1101110010101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1101110010110000000) && ({row_reg, col_reg}<19'b1101110010110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101110010110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1101110010110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1101110010110011010) && ({row_reg, col_reg}<19'b1101110100011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1101110100011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1101110100011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1101110100011101010) && ({row_reg, col_reg}<19'b1101110100011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101110100011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1101110100011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101110100011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1101110100011101111) && ({row_reg, col_reg}<19'b1101110100100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101110100100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1101110100100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1101110100100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1101110100100000100) && ({row_reg, col_reg}<19'b1101110100101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1101110100101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1101110100101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1101110100110000000) && ({row_reg, col_reg}<19'b1101110100110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101110100110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1101110100110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1101110100110011010) && ({row_reg, col_reg}<19'b1101110110011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1101110110011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1101110110011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1101110110011101010) && ({row_reg, col_reg}<19'b1101110110011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101110110011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1101110110011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101110110011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1101110110011101111) && ({row_reg, col_reg}<19'b1101110110100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101110110100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1101110110100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1101110110100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1101110110100000100) && ({row_reg, col_reg}<19'b1101110110101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1101110110101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1101110110101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1101110110110000000) && ({row_reg, col_reg}<19'b1101110110110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101110110110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1101110110110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1101110110110011010) && ({row_reg, col_reg}<19'b1101111000011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1101111000011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1101111000011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1101111000011101010) && ({row_reg, col_reg}<19'b1101111000011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101111000011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1101111000011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101111000011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1101111000011101111) && ({row_reg, col_reg}<19'b1101111000100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101111000100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1101111000100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1101111000100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1101111000100000100) && ({row_reg, col_reg}<19'b1101111000101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1101111000101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1101111000101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1101111000110000000) && ({row_reg, col_reg}<19'b1101111000110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101111000110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1101111000110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1101111000110011010) && ({row_reg, col_reg}<19'b1101111010011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1101111010011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1101111010011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1101111010011101010) && ({row_reg, col_reg}<19'b1101111010011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101111010011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1101111010011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101111010011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1101111010011101111) && ({row_reg, col_reg}<19'b1101111010100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101111010100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1101111010100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1101111010100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1101111010100000100) && ({row_reg, col_reg}<19'b1101111010101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1101111010101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1101111010101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1101111010110000000) && ({row_reg, col_reg}<19'b1101111010110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101111010110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1101111010110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1101111010110011010) && ({row_reg, col_reg}<19'b1101111100011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1101111100011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1101111100011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1101111100011101010) && ({row_reg, col_reg}<19'b1101111100011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101111100011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1101111100011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101111100011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1101111100011101111) && ({row_reg, col_reg}<19'b1101111100100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101111100100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1101111100100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1101111100100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1101111100100000100) && ({row_reg, col_reg}<19'b1101111100101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1101111100101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1101111100101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1101111100110000000) && ({row_reg, col_reg}<19'b1101111100110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101111100110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1101111100110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1101111100110011010) && ({row_reg, col_reg}<19'b1101111110011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1101111110011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1101111110011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1101111110011101010) && ({row_reg, col_reg}<19'b1101111110011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101111110011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1101111110011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101111110011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1101111110011101111) && ({row_reg, col_reg}<19'b1101111110100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101111110100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1101111110100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1101111110100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1101111110100000100) && ({row_reg, col_reg}<19'b1101111110101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1101111110101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1101111110101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1101111110110000000) && ({row_reg, col_reg}<19'b1101111110110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101111110110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1101111110110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1101111110110011010) && ({row_reg, col_reg}<19'b1110000000011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1110000000011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1110000000011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1110000000011101010) && ({row_reg, col_reg}<19'b1110000000011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110000000011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1110000000011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110000000011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1110000000011101111) && ({row_reg, col_reg}<19'b1110000000100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110000000100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1110000000100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1110000000100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1110000000100000100) && ({row_reg, col_reg}<19'b1110000000101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1110000000101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1110000000101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1110000000110000000) && ({row_reg, col_reg}<19'b1110000000110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110000000110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1110000000110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1110000000110011010) && ({row_reg, col_reg}<19'b1110000010011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1110000010011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1110000010011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1110000010011101010) && ({row_reg, col_reg}<19'b1110000010011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110000010011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1110000010011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110000010011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1110000010011101111) && ({row_reg, col_reg}<19'b1110000010100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110000010100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1110000010100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1110000010100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1110000010100000100) && ({row_reg, col_reg}<19'b1110000010101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1110000010101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1110000010101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1110000010110000000) && ({row_reg, col_reg}<19'b1110000010110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110000010110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1110000010110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1110000010110011010) && ({row_reg, col_reg}<19'b1110000100011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1110000100011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1110000100011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1110000100011101010) && ({row_reg, col_reg}<19'b1110000100011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110000100011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1110000100011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110000100011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1110000100011101111) && ({row_reg, col_reg}<19'b1110000100100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110000100100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1110000100100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1110000100100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1110000100100000100) && ({row_reg, col_reg}<19'b1110000100101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1110000100101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1110000100101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1110000100110000000) && ({row_reg, col_reg}<19'b1110000100110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110000100110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1110000100110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1110000100110011010) && ({row_reg, col_reg}<19'b1110000110011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1110000110011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1110000110011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1110000110011101010) && ({row_reg, col_reg}<19'b1110000110011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110000110011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1110000110011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110000110011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1110000110011101111) && ({row_reg, col_reg}<19'b1110000110100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110000110100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1110000110100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1110000110100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1110000110100000100) && ({row_reg, col_reg}<19'b1110000110101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1110000110101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1110000110101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1110000110110000000) && ({row_reg, col_reg}<19'b1110000110110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110000110110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1110000110110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1110000110110011010) && ({row_reg, col_reg}<19'b1110001000011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1110001000011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1110001000011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1110001000011101010) && ({row_reg, col_reg}<19'b1110001000011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110001000011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1110001000011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110001000011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1110001000011101111) && ({row_reg, col_reg}<19'b1110001000100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110001000100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1110001000100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1110001000100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1110001000100000100) && ({row_reg, col_reg}<19'b1110001000101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1110001000101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1110001000101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1110001000110000000) && ({row_reg, col_reg}<19'b1110001000110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110001000110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1110001000110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1110001000110011010) && ({row_reg, col_reg}<19'b1110001010011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1110001010011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1110001010011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1110001010011101010) && ({row_reg, col_reg}<19'b1110001010011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110001010011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1110001010011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110001010011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1110001010011101111) && ({row_reg, col_reg}<19'b1110001010100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110001010100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1110001010100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1110001010100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1110001010100000100) && ({row_reg, col_reg}<19'b1110001010101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1110001010101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1110001010101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1110001010110000000) && ({row_reg, col_reg}<19'b1110001010110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110001010110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1110001010110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1110001010110011010) && ({row_reg, col_reg}<19'b1110001100011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1110001100011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1110001100011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1110001100011101010) && ({row_reg, col_reg}<19'b1110001100011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110001100011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1110001100011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110001100011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1110001100011101111) && ({row_reg, col_reg}<19'b1110001100100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110001100100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1110001100100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1110001100100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1110001100100000100) && ({row_reg, col_reg}<19'b1110001100101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1110001100101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1110001100101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1110001100110000000) && ({row_reg, col_reg}<19'b1110001100110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110001100110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1110001100110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1110001100110011010) && ({row_reg, col_reg}<19'b1110001110011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1110001110011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1110001110011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1110001110011101010) && ({row_reg, col_reg}<19'b1110001110011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110001110011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1110001110011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110001110011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1110001110011101111) && ({row_reg, col_reg}<19'b1110001110100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110001110100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1110001110100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1110001110100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1110001110100000100) && ({row_reg, col_reg}<19'b1110001110101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1110001110101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1110001110101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1110001110110000000) && ({row_reg, col_reg}<19'b1110001110110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110001110110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1110001110110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1110001110110011010) && ({row_reg, col_reg}<19'b1110010000011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1110010000011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1110010000011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1110010000011101010) && ({row_reg, col_reg}<19'b1110010000011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110010000011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1110010000011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110010000011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1110010000011101111) && ({row_reg, col_reg}<19'b1110010000100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110010000100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1110010000100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1110010000100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1110010000100000100) && ({row_reg, col_reg}<19'b1110010000101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1110010000101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1110010000101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1110010000110000000) && ({row_reg, col_reg}<19'b1110010000110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110010000110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1110010000110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1110010000110011010) && ({row_reg, col_reg}<19'b1110010010011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1110010010011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1110010010011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1110010010011101010) && ({row_reg, col_reg}<19'b1110010010011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110010010011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1110010010011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110010010011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1110010010011101111) && ({row_reg, col_reg}<19'b1110010010100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110010010100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1110010010100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1110010010100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1110010010100000100) && ({row_reg, col_reg}<19'b1110010010101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1110010010101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1110010010101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1110010010110000000) && ({row_reg, col_reg}<19'b1110010010110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110010010110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1110010010110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1110010010110011010) && ({row_reg, col_reg}<19'b1110010100011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1110010100011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1110010100011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1110010100011101010) && ({row_reg, col_reg}<19'b1110010100011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110010100011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1110010100011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110010100011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1110010100011101111) && ({row_reg, col_reg}<19'b1110010100100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110010100100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1110010100100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1110010100100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1110010100100000100) && ({row_reg, col_reg}<19'b1110010100101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1110010100101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1110010100101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1110010100110000000) && ({row_reg, col_reg}<19'b1110010100110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110010100110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1110010100110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1110010100110011010) && ({row_reg, col_reg}<19'b1110010110011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1110010110011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1110010110011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1110010110011101010) && ({row_reg, col_reg}<19'b1110010110011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110010110011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1110010110011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110010110011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1110010110011101111) && ({row_reg, col_reg}<19'b1110010110100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110010110100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1110010110100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1110010110100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1110010110100000100) && ({row_reg, col_reg}<19'b1110010110101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1110010110101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1110010110101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1110010110110000000) && ({row_reg, col_reg}<19'b1110010110110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110010110110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1110010110110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1110010110110011010) && ({row_reg, col_reg}<19'b1110011000011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1110011000011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1110011000011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1110011000011101010) && ({row_reg, col_reg}<19'b1110011000011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110011000011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1110011000011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110011000011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1110011000011101111) && ({row_reg, col_reg}<19'b1110011000100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110011000100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1110011000100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1110011000100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1110011000100000100) && ({row_reg, col_reg}<19'b1110011000101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1110011000101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1110011000101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1110011000110000000) && ({row_reg, col_reg}<19'b1110011000110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110011000110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1110011000110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1110011000110011010) && ({row_reg, col_reg}<19'b1110011010011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1110011010011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1110011010011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1110011010011101010) && ({row_reg, col_reg}<19'b1110011010011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110011010011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1110011010011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110011010011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1110011010011101111) && ({row_reg, col_reg}<19'b1110011010100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110011010100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1110011010100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1110011010100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1110011010100000100) && ({row_reg, col_reg}<19'b1110011010101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1110011010101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1110011010101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1110011010110000000) && ({row_reg, col_reg}<19'b1110011010110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110011010110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1110011010110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1110011010110011010) && ({row_reg, col_reg}<19'b1110011100011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1110011100011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1110011100011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1110011100011101010) && ({row_reg, col_reg}<19'b1110011100011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110011100011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1110011100011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110011100011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1110011100011101111) && ({row_reg, col_reg}<19'b1110011100100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110011100100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1110011100100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1110011100100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1110011100100000100) && ({row_reg, col_reg}<19'b1110011100101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1110011100101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1110011100101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1110011100110000000) && ({row_reg, col_reg}<19'b1110011100110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110011100110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1110011100110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1110011100110011010) && ({row_reg, col_reg}<19'b1110011110011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1110011110011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1110011110011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1110011110011101010) && ({row_reg, col_reg}<19'b1110011110011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110011110011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1110011110011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110011110011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1110011110011101111) && ({row_reg, col_reg}<19'b1110011110100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110011110100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1110011110100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1110011110100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1110011110100000100) && ({row_reg, col_reg}<19'b1110011110101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1110011110101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1110011110101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1110011110110000000) && ({row_reg, col_reg}<19'b1110011110110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110011110110011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1110011110110011001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1110011110110011010) && ({row_reg, col_reg}<19'b1110100000011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1110100000011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1110100000011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1110100000011101010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110100000011101011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1110100000011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b1110100000011101101) && ({row_reg, col_reg}<19'b1110100000011110000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1110100000011110000) && ({row_reg, col_reg}<19'b1110100000100000000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b1110100000100000000) && ({row_reg, col_reg}<19'b1110100000100000010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1110100000100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1110100000100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1110100000100000100) && ({row_reg, col_reg}<19'b1110100000101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1110100000101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1110100000101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1110100000110000000) && ({row_reg, col_reg}<19'b1110100000110010000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110100000110010000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1110100000110010001) && ({row_reg, col_reg}<19'b1110100000110010011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b1110100000110010011) && ({row_reg, col_reg}<19'b1110100000110010101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1110100000110010101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110100000110010110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1110100000110010111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110100000110011000)) color_data = 12'b101010101010;

		if(({row_reg, col_reg}>=19'b1110100000110011001) && ({row_reg, col_reg}<19'b1110100010011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1110100010011101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1110100010011101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1110100010011101010) && ({row_reg, col_reg}<19'b1110100010100000010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110100010100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1110100010100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1110100010100000100) && ({row_reg, col_reg}<19'b1110100010101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1110100010101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1110100010101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1110100010110000000) && ({row_reg, col_reg}<19'b1110100010110010000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110100010110010000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1110100010110010001) && ({row_reg, col_reg}<19'b1110100010110011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110100010110011000)) color_data = 12'b101010101010;

		if(({row_reg, col_reg}>=19'b1110100010110011001) && ({row_reg, col_reg}<19'b1110100100011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1110100100011101000)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1110100100011101001) && ({row_reg, col_reg}<19'b1110100100011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1110100100011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110100100011101101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1110100100011101110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110100100011101111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1110100100011110000) && ({row_reg, col_reg}<19'b1110100100100000010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110100100100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1110100100100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1110100100100000100) && ({row_reg, col_reg}<19'b1110100100101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1110100100101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1110100100101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1110100100110000000) && ({row_reg, col_reg}<19'b1110100100110010010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110100100110010010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1110100100110010011) && ({row_reg, col_reg}<19'b1110100100110010111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110100100110010111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1110100100110011000)) color_data = 12'b101010101010;

		if(({row_reg, col_reg}>=19'b1110100100110011001) && ({row_reg, col_reg}<19'b1110100110011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1110100110011101000)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1110100110011101001) && ({row_reg, col_reg}<19'b1110100110011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1110100110011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110100110011101101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1110100110011101110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110100110011101111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1110100110011110000) && ({row_reg, col_reg}<19'b1110100110100000000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b1110100110100000000) && ({row_reg, col_reg}<19'b1110100110100000010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1110100110100000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1110100110100000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1110100110100000100) && ({row_reg, col_reg}<19'b1110100110101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1110100110101111110)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1110100110101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1110100110110000000) && ({row_reg, col_reg}<19'b1110100110110010010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110100110110010010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1110100110110010011) && ({row_reg, col_reg}<19'b1110100110110010101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110100110110010101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1110100110110010110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110100110110010111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1110100110110011000)) color_data = 12'b101010101010;

		if(({row_reg, col_reg}>=19'b1110100110110011001) && ({row_reg, col_reg}<19'b1110101000011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1110101000011101000)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b1110101000011101001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1110101000011101010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110101000011101011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1110101000011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110101000011101101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1110101000011101110) && ({row_reg, col_reg}<19'b1110101000100000000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b1110101000100000000) && ({row_reg, col_reg}<19'b1110101000100000010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1110101000100000010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1110101000100000011)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=19'b1110101000100000100) && ({row_reg, col_reg}<19'b1110101000101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1110101000101111110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b1110101000101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1110101000110000000) && ({row_reg, col_reg}<19'b1110101000110010010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110101000110010010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1110101000110010011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b1110101000110010100) && ({row_reg, col_reg}<19'b1110101000110010110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1110101000110010110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110101000110010111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1110101000110011000)) color_data = 12'b101110111011;

		if(({row_reg, col_reg}>=19'b1110101000110011001) && ({row_reg, col_reg}<19'b1110101010011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1110101010011101000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b1110101010011101001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=19'b1110101010011101010) && ({row_reg, col_reg}<19'b1110101010011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1110101010011101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110101010011101101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1110101010011101110) && ({row_reg, col_reg}<19'b1110101010100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110101010100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1110101010100000010)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=19'b1110101010100000011) && ({row_reg, col_reg}<19'b1110101010101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1110101010101111110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b1110101010101111111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=19'b1110101010110000000) && ({row_reg, col_reg}<19'b1110101010110010000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110101010110010000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1110101010110010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110101010110010010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1110101010110010011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b1110101010110010100) && ({row_reg, col_reg}<19'b1110101010110010110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1110101010110010110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110101010110010111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1110101010110011000)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=19'b1110101010110011001) && ({row_reg, col_reg}<19'b1110101100011101001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1110101100011101001)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=19'b1110101100011101010) && ({row_reg, col_reg}<19'b1110101100011110000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1110101100011110000) && ({row_reg, col_reg}<19'b1110101100100000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110101100100000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1110101100100000010)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=19'b1110101100100000011) && ({row_reg, col_reg}<19'b1110101100101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1110101100101111110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b1110101100101111111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=19'b1110101100110000000) && ({row_reg, col_reg}<19'b1110101100110000011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1110101100110000011) && ({row_reg, col_reg}<19'b1110101100110010000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110101100110010000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1110101100110010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110101100110010010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1110101100110010011) && ({row_reg, col_reg}<19'b1110101100110010111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110101100110010111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1110101100110011000)) color_data = 12'b110111011101;

		if(({row_reg, col_reg}>=19'b1110101100110011001) && ({row_reg, col_reg}<19'b1110101110011101001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1110101110011101001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1110101110011101010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1110101110011101011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110101110011101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1110101110011101101) && ({row_reg, col_reg}<19'b1110101110100000000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110101110100000000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1110101110100000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1110101110100000010)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1110101110100000011) && ({row_reg, col_reg}<19'b1110101110101111111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1110101110101111111)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=19'b1110101110110000000) && ({row_reg, col_reg}<19'b1110101110110000011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1110101110110000011) && ({row_reg, col_reg}<19'b1110101110110010010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110101110110010010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1110101110110010011) && ({row_reg, col_reg}<19'b1110101110110010110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110101110110010110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1110101110110010111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1110101110110011000)) color_data = 12'b110111011101;

		if(({row_reg, col_reg}>=19'b1110101110110011001) && ({row_reg, col_reg}<19'b1110110000011101001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1110110000011101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b1110110000011101010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=19'b1110110000011101011) && ({row_reg, col_reg}<19'b1110110000011101101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1110110000011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110110000011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1110110000011101111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110110000011110000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1110110000011110001) && ({row_reg, col_reg}<19'b1110110000011110100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b1110110000011110100) && ({row_reg, col_reg}<19'b1110110000011110111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1110110000011110111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110110000011111000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1110110000011111001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110110000011111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1110110000011111011) && ({row_reg, col_reg}<19'b1110110000011111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110110000011111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1110110000011111111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110110000100000000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1110110000100000001)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1110110000100000010)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=19'b1110110000100000011) && ({row_reg, col_reg}<19'b1110110000101111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1110110000101111110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b1110110000101111111)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b1110110000110000000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1110110000110000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b1110110000110000010) && ({row_reg, col_reg}<19'b1110110000110000100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1110110000110000100) && ({row_reg, col_reg}<19'b1110110000110000110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110110000110000110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1110110000110000111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b1110110000110001000) && ({row_reg, col_reg}<19'b1110110000110001010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1110110000110001010) && ({row_reg, col_reg}<19'b1110110000110001111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b1110110000110001111) && ({row_reg, col_reg}<19'b1110110000110010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1110110000110010001) && ({row_reg, col_reg}<19'b1110110000110010100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110110000110010100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1110110000110010101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110110000110010110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1110110000110010111)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=19'b1110110000110011000) && ({row_reg, col_reg}<19'b1110110010011101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1110110010011101000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b1110110010011101001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1110110010011101010)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1110110010011101011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1110110010011101100) && ({row_reg, col_reg}<19'b1110110010011110001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b1110110010011110001) && ({row_reg, col_reg}<19'b1110110010011110011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1110110010011110011) && ({row_reg, col_reg}<19'b1110110010011111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b1110110010011111100) && ({row_reg, col_reg}<19'b1110110010011111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1110110010011111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110110010011111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1110110010100000000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1110110010100000001)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1110110010100000010) && ({row_reg, col_reg}<19'b1110110010101111111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1110110010101111111)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b1110110010110000000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1110110010110000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1110110010110000010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b1110110010110000011) && ({row_reg, col_reg}<19'b1110110010110000101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1110110010110000101) && ({row_reg, col_reg}<19'b1110110010110000111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110110010110000111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1110110010110001000) && ({row_reg, col_reg}<19'b1110110010110001011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b1110110010110001011) && ({row_reg, col_reg}<19'b1110110010110001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1110110010110001110) && ({row_reg, col_reg}<19'b1110110010110010000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b1110110010110010000) && ({row_reg, col_reg}<19'b1110110010110010110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1110110010110010110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1110110010110010111)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1110110010110011000) && ({row_reg, col_reg}<19'b1110110100011101010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1110110100011101010)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b1110110100011101011)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=19'b1110110100011101100) && ({row_reg, col_reg}<19'b1110110100011110010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1110110100011110010) && ({row_reg, col_reg}<19'b1110110100011110100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b1110110100011110100) && ({row_reg, col_reg}<19'b1110110100011111000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1110110100011111000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b1110110100011111001) && ({row_reg, col_reg}<19'b1110110100011111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1110110100011111011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b1110110100011111100) && ({row_reg, col_reg}<19'b1110110100100000000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1110110100100000000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1110110100100000001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=19'b1110110100100000010) && ({row_reg, col_reg}<19'b1110110100110000000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1110110100110000000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b1110110100110000001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=19'b1110110100110000010) && ({row_reg, col_reg}<19'b1110110100110000100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110110100110000100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1110110100110000101) && ({row_reg, col_reg}<19'b1110110100110000111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b1110110100110000111) && ({row_reg, col_reg}<19'b1110110100110001001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1110110100110001001) && ({row_reg, col_reg}<19'b1110110100110001111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110110100110001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1110110100110010000) && ({row_reg, col_reg}<19'b1110110100110010011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110110100110010011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1110110100110010100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110110100110010101)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1110110100110010110)) color_data = 12'b110111011101;

		if(({row_reg, col_reg}>=19'b1110110100110010111) && ({row_reg, col_reg}<19'b1110110110011101011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1110110110011101011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b1110110110011101100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1110110110011101101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1110110110011101110) && ({row_reg, col_reg}<19'b1110110110011111011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b1110110110011111011) && ({row_reg, col_reg}<19'b1110110110011111101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1110110110011111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110110110011111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1110110110011111111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1110110110100000000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=19'b1110110110100000001) && ({row_reg, col_reg}<19'b1110110110110000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1110110110110000001)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b1110110110110000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=19'b1110110110110000011) && ({row_reg, col_reg}<19'b1110110110110000110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110110110110000110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1110110110110000111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b1110110110110001000) && ({row_reg, col_reg}<19'b1110110110110001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1110110110110001110) && ({row_reg, col_reg}<19'b1110110110110010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110110110110010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1110110110110010010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b1110110110110010011) && ({row_reg, col_reg}<19'b1110110110110010101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1110110110110010101)) color_data = 12'b101110111011;

		if(({row_reg, col_reg}>=19'b1110110110110010110) && ({row_reg, col_reg}<19'b1110111000011101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1110111000011101100)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b1110111000011101101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1110111000011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1110111000011101111) && ({row_reg, col_reg}<19'b1110111000011110001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b1110111000011110001) && ({row_reg, col_reg}<19'b1110111000011110100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1110111000011110100) && ({row_reg, col_reg}<19'b1110111000011110111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b1110111000011110111) && ({row_reg, col_reg}<19'b1110111000011111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1110111000011111001) && ({row_reg, col_reg}<19'b1110111000011111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110111000011111101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1110111000011111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1110111000011111111)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=19'b1110111000100000000) && ({row_reg, col_reg}<19'b1110111000110000010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1110111000110000010)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1110111000110000011)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1110111000110000100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1110111000110000101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b1110111000110000110) && ({row_reg, col_reg}<19'b1110111000110001000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1110111000110001000) && ({row_reg, col_reg}<19'b1110111000110010000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110111000110010000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1110111000110010001) && ({row_reg, col_reg}<19'b1110111000110010011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110111000110010011)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1110111000110010100)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1110111000110010101)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1110111000110010110) && ({row_reg, col_reg}<19'b1110111010011101010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1110111010011101010)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=19'b1110111010011101011) && ({row_reg, col_reg}<19'b1110111010011101101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1110111010011101101)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b1110111010011101110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1110111010011101111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1110111010011110000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1110111010011110001) && ({row_reg, col_reg}<19'b1110111010011110100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110111010011110100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1110111010011110101) && ({row_reg, col_reg}<19'b1110111010011110111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110111010011110111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1110111010011111000) && ({row_reg, col_reg}<19'b1110111010011111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110111010011111100)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1110111010011111101)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=19'b1110111010011111110) && ({row_reg, col_reg}<19'b1110111010110000011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1110111010110000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b1110111010110000100)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1110111010110000101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1110111010110000110) && ({row_reg, col_reg}<19'b1110111010110001011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b1110111010110001011) && ({row_reg, col_reg}<19'b1110111010110010010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1110111010110010010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1110111010110010011)) color_data = 12'b110111011101;

		if(({row_reg, col_reg}>=19'b1110111010110010100) && ({row_reg, col_reg}<19'b1110111100011101111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1110111100011101111)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1110111100011110000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1110111100011110001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=19'b1110111100011110010) && ({row_reg, col_reg}<19'b1110111100011110101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1110111100011110101) && ({row_reg, col_reg}<19'b1110111100011110111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b1110111100011110111) && ({row_reg, col_reg}<19'b1110111100011111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1110111100011111010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1110111100011111011)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1110111100011111100)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1110111100011111101) && ({row_reg, col_reg}<19'b1110111100110000100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1110111100110000100)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b1110111100110000101)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1110111100110000110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=19'b1110111100110000111) && ({row_reg, col_reg}<19'b1110111100110001011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1110111100110001011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b1110111100110001100) && ({row_reg, col_reg}<19'b1110111100110010000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1110111100110010000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1110111100110010001)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1110111100110010010)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1110111100110010011) && ({row_reg, col_reg}<19'b1110111110011110000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1110111110011110000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b1110111110011110001)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b1110111110011110010)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1110111110011110011)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1110111110011110100)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=19'b1110111110011110101) && ({row_reg, col_reg}<19'b1110111110011110111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1110111110011110111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1110111110011111000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1110111110011111001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1110111110011111010)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b1110111110011111011)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=19'b1110111110011111100) && ({row_reg, col_reg}<19'b1110111110110000110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1110111110110000110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b1110111110110000111)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1110111110110001000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1110111110110001001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1110111110110001010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=19'b1110111110110001011) && ({row_reg, col_reg}<19'b1110111110110001101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1110111110110001101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1110111110110001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1110111110110001111)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1110111110110010000)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b1110111110110010001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1110111110110010010) && ({row_reg, col_reg}<=19'b1110111111001111111)) color_data = 12'b111111111111;
	end
endmodule