module tictactoeboard_rom
	(
		input wire clk,
		input wire [8:0] row,
		input wire [9:0] col,
		output reg [11:0] color_data
	);

	(* rom_style = "block" *)

	//signal declaration
	reg [8:0] row_reg;
	reg [9:0] col_reg;

	always @(posedge clk)
		begin
		row_reg <= row;
		col_reg <= col;
		end

	always @(*) begin
		if(({row_reg, col_reg}>=19'b0000000000000000000) && ({row_reg, col_reg}<19'b0000000000101000000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0000000000101000000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0000000000101000001)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0000000000101000010)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0000000000101000011)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0000000000101000100)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0000000000101000101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0000000000101000110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0000000000101000111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0000000000101001000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0000000000101001001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0000000000101001010)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0000000000101001011)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=19'b0000000000101001100) && ({row_reg, col_reg}<19'b0000000000111010110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=19'b0000000000111010110) && ({row_reg, col_reg}<19'b0000000000111011000)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0000000000111011000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0000000000111011001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0000000000111011010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0000000000111011011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0000000000111011100)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0000000000111011101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0000000000111011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0000000000111011111)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0000000000111100000)) color_data = 12'b110111011101;

		if(({row_reg, col_reg}>=19'b0000000000111100001) && ({row_reg, col_reg}<19'b0000000010100111110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0000000010100111110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0000000010100111111)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0000000010101000000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0000000010101000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=19'b0000000010101000010) && ({row_reg, col_reg}<19'b0000000010101000110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000000010101000110) && ({row_reg, col_reg}<19'b0000000010101001000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0000000010101001000) && ({row_reg, col_reg}<19'b0000000010101001010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0000000010101001010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0000000010101001011)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0000000010101001100)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=19'b0000000010101001101) && ({row_reg, col_reg}<19'b0000000010111010100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0000000010111010100)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0000000010111010101)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0000000010111010110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=19'b0000000010111010111) && ({row_reg, col_reg}<19'b0000000010111011010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000000010111011010) && ({row_reg, col_reg}<19'b0000000010111011100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0000000010111011100) && ({row_reg, col_reg}<19'b0000000010111100000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0000000010111100000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0000000010111100001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0000000010111100010)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0000000010111100011) && ({row_reg, col_reg}<19'b0000000100100111101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0000000100100111101)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0000000100100111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0000000100100111111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0000000100101000000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000000100101000001) && ({row_reg, col_reg}<19'b0000000100101000111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000000100101000111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0000000100101001000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000000100101001001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000000100101001010) && ({row_reg, col_reg}<19'b0000000100101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000000100101001100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0000000100101001101)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0000000100101001110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=19'b0000000100101001111) && ({row_reg, col_reg}<19'b0000000100111010011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0000000100111010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0000000100111010100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=19'b0000000100111010101) && ({row_reg, col_reg}<19'b0000000100111010111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0000000100111010111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000000100111011000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0000000100111011001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0000000100111011010) && ({row_reg, col_reg}<19'b0000000100111011101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000000100111011101) && ({row_reg, col_reg}<19'b0000000100111011111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0000000100111011111) && ({row_reg, col_reg}<19'b0000000100111100010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0000000100111100010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0000000100111100011)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0000000100111100100)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0000000100111100101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0000000100111100110)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0000000100111100111) && ({row_reg, col_reg}<19'b0000000110100111100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0000000110100111100)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0000000110100111101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=19'b0000000110100111110) && ({row_reg, col_reg}<19'b0000000110101000000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0000000110101000000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0000000110101000001) && ({row_reg, col_reg}<19'b0000000110101001011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0000000110101001011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0000000110101001100) && ({row_reg, col_reg}<19'b0000000110101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0000000110101001110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0000000110101001111)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=19'b0000000110101010000) && ({row_reg, col_reg}<19'b0000000110111010010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0000000110111010010)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0000000110111010011)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0000000110111010100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000000110111010101) && ({row_reg, col_reg}<19'b0000000110111010111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000000110111010111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000000110111011000) && ({row_reg, col_reg}<19'b0000000110111100010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000000110111100010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0000000110111100011)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0000000110111100100)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0000000110111100101)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0000000110111100110) && ({row_reg, col_reg}<19'b0000001000100111011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0000001000100111011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0000001000100111100)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0000001000100111101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0000001000100111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000001000100111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000001000101000000) && ({row_reg, col_reg}<19'b0000001000101001010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0000001000101001010) && ({row_reg, col_reg}<19'b0000001000101001101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0000001000101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000001000101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0000001000101001111)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0000001000101010000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=19'b0000001000101010001) && ({row_reg, col_reg}<19'b0000001000111010001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0000001000111010001)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0000001000111010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0000001000111010011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0000001000111010100) && ({row_reg, col_reg}<19'b0000001000111010110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000001000111010110) && ({row_reg, col_reg}<19'b0000001000111011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0000001000111011000) && ({row_reg, col_reg}<19'b0000001000111011110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000001000111011110) && ({row_reg, col_reg}<19'b0000001000111100011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0000001000111100011) && ({row_reg, col_reg}<19'b0000001000111100101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0000001000111100101)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=19'b0000001000111100110) && ({row_reg, col_reg}<19'b0000001010100111010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0000001010100111010)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0000001010100111011)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=19'b0000001010100111100) && ({row_reg, col_reg}<19'b0000001010100111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000001010100111111) && ({row_reg, col_reg}<19'b0000001010101000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0000001010101000001) && ({row_reg, col_reg}<19'b0000001010101000100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000001010101000100) && ({row_reg, col_reg}<19'b0000001010101000110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0000001010101000110) && ({row_reg, col_reg}<19'b0000001010101001011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000001010101001011) && ({row_reg, col_reg}<19'b0000001010101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0000001010101001101) && ({row_reg, col_reg}<19'b0000001010101010000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0000001010101010000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0000001010101010001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=19'b0000001010101010010) && ({row_reg, col_reg}<19'b0000001010111010000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0000001010111010000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0000001010111010001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0000001010111010010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000001010111010011) && ({row_reg, col_reg}<19'b0000001010111010111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0000001010111010111) && ({row_reg, col_reg}<19'b0000001010111011010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000001010111011010) && ({row_reg, col_reg}<19'b0000001010111100000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000001010111100000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000001010111100001) && ({row_reg, col_reg}<19'b0000001010111100011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000001010111100011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0000001010111100100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000001010111100101)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0000001010111100110)) color_data = 12'b110111011101;

		if(({row_reg, col_reg}>=19'b0000001010111100111) && ({row_reg, col_reg}<19'b0000001100100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0000001100100111000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0000001100100111001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0000001100100111010)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0000001100100111011)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=19'b0000001100100111100) && ({row_reg, col_reg}<19'b0000001100100111111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000001100100111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000001100101000000) && ({row_reg, col_reg}<19'b0000001100101000101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000001100101000101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000001100101000110) && ({row_reg, col_reg}<19'b0000001100101001000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000001100101001000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000001100101001001) && ({row_reg, col_reg}<19'b0000001100101001011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0000001100101001011) && ({row_reg, col_reg}<19'b0000001100101001101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000001100101001101) && ({row_reg, col_reg}<19'b0000001100101001111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000001100101001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0000001100101010000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0000001100101010001)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0000001100101010010) && ({row_reg, col_reg}<19'b0000001100111001111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0000001100111001111)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0000001100111010000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0000001100111010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000001100111010010) && ({row_reg, col_reg}<19'b0000001100111010101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000001100111010101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0000001100111010110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000001100111010111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000001100111011000) && ({row_reg, col_reg}<19'b0000001100111011010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0000001100111011010) && ({row_reg, col_reg}<19'b0000001100111011110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000001100111011110) && ({row_reg, col_reg}<19'b0000001100111100001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0000001100111100001) && ({row_reg, col_reg}<19'b0000001100111100011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000001100111100011) && ({row_reg, col_reg}<19'b0000001100111100101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000001100111100101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0000001100111100110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0000001100111100111)) color_data = 12'b110111011101;

		if(({row_reg, col_reg}>=19'b0000001100111101000) && ({row_reg, col_reg}<19'b0000001110100111001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0000001110100111001)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0000001110100111010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0000001110100111011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0000001110100111100) && ({row_reg, col_reg}<19'b0000001110100111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000001110100111111) && ({row_reg, col_reg}<19'b0000001110101000111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000001110101000111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000001110101001000) && ({row_reg, col_reg}<19'b0000001110101001010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0000001110101001010) && ({row_reg, col_reg}<19'b0000001110101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000001110101001100) && ({row_reg, col_reg}<19'b0000001110101001110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000001110101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000001110101001111) && ({row_reg, col_reg}<19'b0000001110101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000001110101010001)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0000001110101010010)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=19'b0000001110101010011) && ({row_reg, col_reg}<19'b0000001110111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0000001110111001110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0000001110111001111)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0000001110111010000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0000001110111010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000001110111010010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000001110111010011) && ({row_reg, col_reg}<19'b0000001110111010101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000001110111010101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000001110111010110) && ({row_reg, col_reg}<19'b0000001110111011001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0000001110111011001) && ({row_reg, col_reg}<19'b0000001110111011011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000001110111011011) && ({row_reg, col_reg}<19'b0000001110111100000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000001110111100000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000001110111100001) && ({row_reg, col_reg}<19'b0000001110111100100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000001110111100100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0000001110111100101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000001110111100110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0000001110111100111)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=19'b0000001110111101000) && ({row_reg, col_reg}<19'b0000010000100111001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0000010000100111001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0000010000100111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0000010000100111011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000010000100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0000010000100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000010000100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000010000100111111) && ({row_reg, col_reg}<19'b0000010000101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000010000101010001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0000010000101010010)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0000010000101010011) && ({row_reg, col_reg}<19'b0000010000111001111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0000010000111001111)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=19'b0000010000111010000) && ({row_reg, col_reg}<19'b0000010000111010011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000010000111010011) && ({row_reg, col_reg}<19'b0000010000111100010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000010000111100010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000010000111100011) && ({row_reg, col_reg}<19'b0000010000111100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000010000111100110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0000010000111100111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0000010000111101000)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0000010000111101001) && ({row_reg, col_reg}<19'b0000010010100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0000010010100111000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0000010010100111001)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0000010010100111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0000010010100111011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000010010100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000010010100111101) && ({row_reg, col_reg}<19'b0000010010101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000010010101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0000010010101010010)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=19'b0000010010101010011) && ({row_reg, col_reg}<19'b0000010010111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0000010010111001110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0000010010111001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=19'b0000010010111010000) && ({row_reg, col_reg}<19'b0000010010111100000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000010010111100000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0000010010111100001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000010010111100010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000010010111100011) && ({row_reg, col_reg}<19'b0000010010111100111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000010010111100111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0000010010111101000)) color_data = 12'b110111011101;

		if(({row_reg, col_reg}>=19'b0000010010111101001) && ({row_reg, col_reg}<19'b0000010100100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0000010100100111000)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0000010100100111001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0000010100100111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0000010100100111011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000010100100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000010100100111101) && ({row_reg, col_reg}<19'b0000010100100111111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000010100100111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000010100101000000) && ({row_reg, col_reg}<19'b0000010100101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000010100101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0000010100101010010)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=19'b0000010100101010011) && ({row_reg, col_reg}<19'b0000010100111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0000010100111001110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0000010100111001111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=19'b0000010100111010000) && ({row_reg, col_reg}<19'b0000010100111100000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000010100111100000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0000010100111100001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000010100111100010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0000010100111100011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0000010100111100100) && ({row_reg, col_reg}<19'b0000010100111100110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0000010100111100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000010100111100111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0000010100111101000)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=19'b0000010100111101001) && ({row_reg, col_reg}<19'b0000010110100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0000010110100111000)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0000010110100111001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=19'b0000010110100111010) && ({row_reg, col_reg}<19'b0000010110100111101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000010110100111101) && ({row_reg, col_reg}<19'b0000010110100111111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000010110100111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000010110101000000) && ({row_reg, col_reg}<19'b0000010110101010000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0000010110101010000) && ({row_reg, col_reg}<19'b0000010110101010010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0000010110101010010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0000010110101010011)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=19'b0000010110101010100) && ({row_reg, col_reg}<19'b0000010110111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0000010110111001110)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0000010110111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000010110111010000) && ({row_reg, col_reg}<19'b0000010110111100010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000010110111100010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0000010110111100011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0000010110111100100) && ({row_reg, col_reg}<19'b0000010110111100110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0000010110111100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000010110111100111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0000010110111101000)) color_data = 12'b101110111011;

		if(({row_reg, col_reg}>=19'b0000010110111101001) && ({row_reg, col_reg}<19'b0000011000100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0000011000100111000)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0000011000100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0000011000100111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000011000100111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000011000100111100) && ({row_reg, col_reg}<19'b0000011000101010000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0000011000101010000) && ({row_reg, col_reg}<19'b0000011000101010010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0000011000101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0000011000101010011)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=19'b0000011000101010100) && ({row_reg, col_reg}<19'b0000011000111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0000011000111001110)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0000011000111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000011000111010000) && ({row_reg, col_reg}<19'b0000011000111100010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000011000111100010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000011000111100011) && ({row_reg, col_reg}<19'b0000011000111100101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0000011000111100101) && ({row_reg, col_reg}<19'b0000011000111101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0000011000111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0000011000111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0000011000111101010) && ({row_reg, col_reg}<19'b0000011010100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0000011010100111000)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0000011010100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000011010100111010) && ({row_reg, col_reg}<19'b0000011010100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000011010100111101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000011010100111110) && ({row_reg, col_reg}<19'b0000011010101010010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000011010101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0000011010101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0000011010101010100) && ({row_reg, col_reg}<19'b0000011010111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0000011010111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0000011010111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000011010111010000) && ({row_reg, col_reg}<19'b0000011010111100001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0000011010111100001) && ({row_reg, col_reg}<19'b0000011010111100011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000011010111100011) && ({row_reg, col_reg}<19'b0000011010111100111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000011010111100111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0000011010111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0000011010111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0000011010111101010) && ({row_reg, col_reg}<19'b0000011100100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0000011100100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0000011100100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000011100100111010) && ({row_reg, col_reg}<19'b0000011100100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0000011100100111100) && ({row_reg, col_reg}<19'b0000011100100111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000011100100111111) && ({row_reg, col_reg}<19'b0000011100101010010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000011100101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0000011100101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0000011100101010100) && ({row_reg, col_reg}<19'b0000011100111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0000011100111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=19'b0000011100111001111) && ({row_reg, col_reg}<19'b0000011100111010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000011100111010001) && ({row_reg, col_reg}<19'b0000011100111100011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000011100111100011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000011100111100100) && ({row_reg, col_reg}<19'b0000011100111100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000011100111100110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0000011100111100111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000011100111101000)) color_data = 12'b101010101010;

		if(({row_reg, col_reg}>=19'b0000011100111101001) && ({row_reg, col_reg}<19'b0000011110100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0000011110100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=19'b0000011110100111001) && ({row_reg, col_reg}<19'b0000011110100111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0000011110100111011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000011110100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000011110100111101) && ({row_reg, col_reg}<19'b0000011110101010010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000011110101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0000011110101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0000011110101010100) && ({row_reg, col_reg}<19'b0000011110111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0000011110111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0000011110111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000011110111010000) && ({row_reg, col_reg}<19'b0000011110111010111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000011110111010111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000011110111011000) && ({row_reg, col_reg}<19'b0000011110111100000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000011110111100000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000011110111100001) && ({row_reg, col_reg}<19'b0000011110111100011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0000011110111100011) && ({row_reg, col_reg}<19'b0000011110111100101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0000011110111100101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000011110111100110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0000011110111100111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000011110111101000)) color_data = 12'b101010101010;

		if(({row_reg, col_reg}>=19'b0000011110111101001) && ({row_reg, col_reg}<19'b0000100000100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0000100000100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0000100000100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000100000100111010) && ({row_reg, col_reg}<19'b0000100000100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000100000100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0000100000100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000100000100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000100000100111111) && ({row_reg, col_reg}<19'b0000100000101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000100000101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0000100000101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0000100000101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0000100000101010100) && ({row_reg, col_reg}<19'b0000100000111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0000100000111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0000100000111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000100000111010000) && ({row_reg, col_reg}<19'b0000100000111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000100000111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0000100000111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0000100000111101010) && ({row_reg, col_reg}<19'b0000100010100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0000100010100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0000100010100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000100010100111010) && ({row_reg, col_reg}<19'b0000100010100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000100010100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0000100010100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000100010100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000100010100111111) && ({row_reg, col_reg}<19'b0000100010101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000100010101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0000100010101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0000100010101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0000100010101010100) && ({row_reg, col_reg}<19'b0000100010111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0000100010111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0000100010111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000100010111010000) && ({row_reg, col_reg}<19'b0000100010111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000100010111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0000100010111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0000100010111101010) && ({row_reg, col_reg}<19'b0000100100100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0000100100100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0000100100100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000100100100111010) && ({row_reg, col_reg}<19'b0000100100100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000100100100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0000100100100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000100100100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000100100100111111) && ({row_reg, col_reg}<19'b0000100100101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000100100101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0000100100101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0000100100101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0000100100101010100) && ({row_reg, col_reg}<19'b0000100100111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0000100100111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0000100100111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000100100111010000) && ({row_reg, col_reg}<19'b0000100100111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000100100111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0000100100111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0000100100111101010) && ({row_reg, col_reg}<19'b0000100110100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0000100110100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0000100110100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000100110100111010) && ({row_reg, col_reg}<19'b0000100110100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000100110100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0000100110100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000100110100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000100110100111111) && ({row_reg, col_reg}<19'b0000100110101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000100110101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0000100110101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0000100110101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0000100110101010100) && ({row_reg, col_reg}<19'b0000100110111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0000100110111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0000100110111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000100110111010000) && ({row_reg, col_reg}<19'b0000100110111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000100110111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0000100110111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0000100110111101010) && ({row_reg, col_reg}<19'b0000101000100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0000101000100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0000101000100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000101000100111010) && ({row_reg, col_reg}<19'b0000101000100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000101000100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0000101000100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000101000100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000101000100111111) && ({row_reg, col_reg}<19'b0000101000101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000101000101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0000101000101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0000101000101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0000101000101010100) && ({row_reg, col_reg}<19'b0000101000111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0000101000111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0000101000111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000101000111010000) && ({row_reg, col_reg}<19'b0000101000111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000101000111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0000101000111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0000101000111101010) && ({row_reg, col_reg}<19'b0000101010100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0000101010100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0000101010100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000101010100111010) && ({row_reg, col_reg}<19'b0000101010100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000101010100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0000101010100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000101010100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000101010100111111) && ({row_reg, col_reg}<19'b0000101010101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000101010101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0000101010101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0000101010101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0000101010101010100) && ({row_reg, col_reg}<19'b0000101010111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0000101010111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0000101010111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000101010111010000) && ({row_reg, col_reg}<19'b0000101010111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000101010111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0000101010111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0000101010111101010) && ({row_reg, col_reg}<19'b0000101100100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0000101100100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0000101100100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000101100100111010) && ({row_reg, col_reg}<19'b0000101100100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000101100100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0000101100100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000101100100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000101100100111111) && ({row_reg, col_reg}<19'b0000101100101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000101100101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0000101100101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0000101100101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0000101100101010100) && ({row_reg, col_reg}<19'b0000101100111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0000101100111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0000101100111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000101100111010000) && ({row_reg, col_reg}<19'b0000101100111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000101100111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0000101100111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0000101100111101010) && ({row_reg, col_reg}<19'b0000101110100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0000101110100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0000101110100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000101110100111010) && ({row_reg, col_reg}<19'b0000101110100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000101110100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0000101110100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000101110100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000101110100111111) && ({row_reg, col_reg}<19'b0000101110101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000101110101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0000101110101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0000101110101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0000101110101010100) && ({row_reg, col_reg}<19'b0000101110111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0000101110111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0000101110111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000101110111010000) && ({row_reg, col_reg}<19'b0000101110111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000101110111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0000101110111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0000101110111101010) && ({row_reg, col_reg}<19'b0000110000100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0000110000100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0000110000100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000110000100111010) && ({row_reg, col_reg}<19'b0000110000100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000110000100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0000110000100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000110000100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000110000100111111) && ({row_reg, col_reg}<19'b0000110000101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000110000101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0000110000101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0000110000101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0000110000101010100) && ({row_reg, col_reg}<19'b0000110000111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0000110000111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0000110000111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000110000111010000) && ({row_reg, col_reg}<19'b0000110000111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000110000111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0000110000111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0000110000111101010) && ({row_reg, col_reg}<19'b0000110010100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0000110010100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0000110010100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000110010100111010) && ({row_reg, col_reg}<19'b0000110010100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000110010100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0000110010100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000110010100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000110010100111111) && ({row_reg, col_reg}<19'b0000110010101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000110010101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0000110010101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0000110010101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0000110010101010100) && ({row_reg, col_reg}<19'b0000110010111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0000110010111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0000110010111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000110010111010000) && ({row_reg, col_reg}<19'b0000110010111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000110010111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0000110010111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0000110010111101010) && ({row_reg, col_reg}<19'b0000110100100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0000110100100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0000110100100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000110100100111010) && ({row_reg, col_reg}<19'b0000110100100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000110100100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0000110100100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000110100100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000110100100111111) && ({row_reg, col_reg}<19'b0000110100101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000110100101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0000110100101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0000110100101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0000110100101010100) && ({row_reg, col_reg}<19'b0000110100111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0000110100111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0000110100111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000110100111010000) && ({row_reg, col_reg}<19'b0000110100111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000110100111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0000110100111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0000110100111101010) && ({row_reg, col_reg}<19'b0000110110100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0000110110100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0000110110100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000110110100111010) && ({row_reg, col_reg}<19'b0000110110100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000110110100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0000110110100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000110110100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000110110100111111) && ({row_reg, col_reg}<19'b0000110110101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000110110101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0000110110101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0000110110101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0000110110101010100) && ({row_reg, col_reg}<19'b0000110110111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0000110110111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0000110110111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000110110111010000) && ({row_reg, col_reg}<19'b0000110110111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000110110111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0000110110111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0000110110111101010) && ({row_reg, col_reg}<19'b0000111000100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0000111000100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0000111000100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000111000100111010) && ({row_reg, col_reg}<19'b0000111000100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000111000100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0000111000100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000111000100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000111000100111111) && ({row_reg, col_reg}<19'b0000111000101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000111000101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0000111000101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0000111000101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0000111000101010100) && ({row_reg, col_reg}<19'b0000111000111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0000111000111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0000111000111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000111000111010000) && ({row_reg, col_reg}<19'b0000111000111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000111000111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0000111000111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0000111000111101010) && ({row_reg, col_reg}<19'b0000111010100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0000111010100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0000111010100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000111010100111010) && ({row_reg, col_reg}<19'b0000111010100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000111010100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0000111010100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000111010100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000111010100111111) && ({row_reg, col_reg}<19'b0000111010101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000111010101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0000111010101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0000111010101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0000111010101010100) && ({row_reg, col_reg}<19'b0000111010111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0000111010111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0000111010111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000111010111010000) && ({row_reg, col_reg}<19'b0000111010111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000111010111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0000111010111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0000111010111101010) && ({row_reg, col_reg}<19'b0000111100100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0000111100100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0000111100100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000111100100111010) && ({row_reg, col_reg}<19'b0000111100100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000111100100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0000111100100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000111100100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000111100100111111) && ({row_reg, col_reg}<19'b0000111100101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000111100101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0000111100101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0000111100101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0000111100101010100) && ({row_reg, col_reg}<19'b0000111100111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0000111100111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0000111100111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000111100111010000) && ({row_reg, col_reg}<19'b0000111100111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000111100111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0000111100111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0000111100111101010) && ({row_reg, col_reg}<19'b0000111110100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0000111110100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0000111110100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000111110100111010) && ({row_reg, col_reg}<19'b0000111110100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000111110100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0000111110100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000111110100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000111110100111111) && ({row_reg, col_reg}<19'b0000111110101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000111110101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0000111110101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0000111110101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0000111110101010100) && ({row_reg, col_reg}<19'b0000111110111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0000111110111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0000111110111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0000111110111010000) && ({row_reg, col_reg}<19'b0000111110111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0000111110111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0000111110111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0000111110111101010) && ({row_reg, col_reg}<19'b0001000000100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0001000000100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0001000000100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0001000000100111010) && ({row_reg, col_reg}<19'b0001000000100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001000000100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0001000000100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001000000100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0001000000100111111) && ({row_reg, col_reg}<19'b0001000000101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001000000101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0001000000101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0001000000101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0001000000101010100) && ({row_reg, col_reg}<19'b0001000000111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0001000000111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0001000000111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0001000000111010000) && ({row_reg, col_reg}<19'b0001000000111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001000000111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0001000000111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0001000000111101010) && ({row_reg, col_reg}<19'b0001000010100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0001000010100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0001000010100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0001000010100111010) && ({row_reg, col_reg}<19'b0001000010100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001000010100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0001000010100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001000010100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0001000010100111111) && ({row_reg, col_reg}<19'b0001000010101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001000010101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0001000010101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0001000010101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0001000010101010100) && ({row_reg, col_reg}<19'b0001000010111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0001000010111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0001000010111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0001000010111010000) && ({row_reg, col_reg}<19'b0001000010111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001000010111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0001000010111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0001000010111101010) && ({row_reg, col_reg}<19'b0001000100100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0001000100100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0001000100100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0001000100100111010) && ({row_reg, col_reg}<19'b0001000100100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001000100100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0001000100100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001000100100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0001000100100111111) && ({row_reg, col_reg}<19'b0001000100101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001000100101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0001000100101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0001000100101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0001000100101010100) && ({row_reg, col_reg}<19'b0001000100111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0001000100111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0001000100111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0001000100111010000) && ({row_reg, col_reg}<19'b0001000100111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001000100111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0001000100111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0001000100111101010) && ({row_reg, col_reg}<19'b0001000110100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0001000110100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0001000110100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0001000110100111010) && ({row_reg, col_reg}<19'b0001000110100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001000110100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0001000110100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001000110100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0001000110100111111) && ({row_reg, col_reg}<19'b0001000110101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001000110101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0001000110101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0001000110101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0001000110101010100) && ({row_reg, col_reg}<19'b0001000110111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0001000110111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0001000110111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0001000110111010000) && ({row_reg, col_reg}<19'b0001000110111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001000110111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0001000110111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0001000110111101010) && ({row_reg, col_reg}<19'b0001001000100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0001001000100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0001001000100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0001001000100111010) && ({row_reg, col_reg}<19'b0001001000100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001001000100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0001001000100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001001000100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0001001000100111111) && ({row_reg, col_reg}<19'b0001001000101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001001000101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0001001000101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0001001000101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0001001000101010100) && ({row_reg, col_reg}<19'b0001001000111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0001001000111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0001001000111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0001001000111010000) && ({row_reg, col_reg}<19'b0001001000111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001001000111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0001001000111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0001001000111101010) && ({row_reg, col_reg}<19'b0001001010100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0001001010100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0001001010100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0001001010100111010) && ({row_reg, col_reg}<19'b0001001010100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001001010100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0001001010100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001001010100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0001001010100111111) && ({row_reg, col_reg}<19'b0001001010101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001001010101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0001001010101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0001001010101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0001001010101010100) && ({row_reg, col_reg}<19'b0001001010111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0001001010111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0001001010111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0001001010111010000) && ({row_reg, col_reg}<19'b0001001010111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001001010111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0001001010111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0001001010111101010) && ({row_reg, col_reg}<19'b0001001100100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0001001100100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0001001100100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0001001100100111010) && ({row_reg, col_reg}<19'b0001001100100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001001100100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0001001100100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001001100100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0001001100100111111) && ({row_reg, col_reg}<19'b0001001100101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001001100101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0001001100101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0001001100101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0001001100101010100) && ({row_reg, col_reg}<19'b0001001100111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0001001100111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0001001100111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0001001100111010000) && ({row_reg, col_reg}<19'b0001001100111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001001100111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0001001100111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0001001100111101010) && ({row_reg, col_reg}<19'b0001001110100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0001001110100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0001001110100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0001001110100111010) && ({row_reg, col_reg}<19'b0001001110100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001001110100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0001001110100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001001110100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0001001110100111111) && ({row_reg, col_reg}<19'b0001001110101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001001110101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0001001110101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0001001110101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0001001110101010100) && ({row_reg, col_reg}<19'b0001001110111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0001001110111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0001001110111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0001001110111010000) && ({row_reg, col_reg}<19'b0001001110111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001001110111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0001001110111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0001001110111101010) && ({row_reg, col_reg}<19'b0001010000100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0001010000100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0001010000100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0001010000100111010) && ({row_reg, col_reg}<19'b0001010000100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001010000100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0001010000100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001010000100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0001010000100111111) && ({row_reg, col_reg}<19'b0001010000101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001010000101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0001010000101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0001010000101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0001010000101010100) && ({row_reg, col_reg}<19'b0001010000111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0001010000111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0001010000111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0001010000111010000) && ({row_reg, col_reg}<19'b0001010000111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001010000111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0001010000111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0001010000111101010) && ({row_reg, col_reg}<19'b0001010010100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0001010010100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0001010010100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0001010010100111010) && ({row_reg, col_reg}<19'b0001010010100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001010010100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0001010010100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001010010100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0001010010100111111) && ({row_reg, col_reg}<19'b0001010010101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001010010101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0001010010101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0001010010101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0001010010101010100) && ({row_reg, col_reg}<19'b0001010010111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0001010010111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0001010010111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0001010010111010000) && ({row_reg, col_reg}<19'b0001010010111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001010010111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0001010010111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0001010010111101010) && ({row_reg, col_reg}<19'b0001010100100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0001010100100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0001010100100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0001010100100111010) && ({row_reg, col_reg}<19'b0001010100100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001010100100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0001010100100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001010100100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0001010100100111111) && ({row_reg, col_reg}<19'b0001010100101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001010100101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0001010100101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0001010100101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0001010100101010100) && ({row_reg, col_reg}<19'b0001010100111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0001010100111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0001010100111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0001010100111010000) && ({row_reg, col_reg}<19'b0001010100111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001010100111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0001010100111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0001010100111101010) && ({row_reg, col_reg}<19'b0001010110100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0001010110100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0001010110100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0001010110100111010) && ({row_reg, col_reg}<19'b0001010110100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001010110100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0001010110100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001010110100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0001010110100111111) && ({row_reg, col_reg}<19'b0001010110101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001010110101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0001010110101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0001010110101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0001010110101010100) && ({row_reg, col_reg}<19'b0001010110111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0001010110111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0001010110111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0001010110111010000) && ({row_reg, col_reg}<19'b0001010110111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001010110111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0001010110111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0001010110111101010) && ({row_reg, col_reg}<19'b0001011000100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0001011000100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0001011000100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0001011000100111010) && ({row_reg, col_reg}<19'b0001011000100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001011000100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0001011000100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001011000100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0001011000100111111) && ({row_reg, col_reg}<19'b0001011000101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001011000101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0001011000101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0001011000101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0001011000101010100) && ({row_reg, col_reg}<19'b0001011000111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0001011000111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0001011000111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0001011000111010000) && ({row_reg, col_reg}<19'b0001011000111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001011000111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0001011000111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0001011000111101010) && ({row_reg, col_reg}<19'b0001011010100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0001011010100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0001011010100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0001011010100111010) && ({row_reg, col_reg}<19'b0001011010100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001011010100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0001011010100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001011010100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0001011010100111111) && ({row_reg, col_reg}<19'b0001011010101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001011010101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0001011010101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0001011010101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0001011010101010100) && ({row_reg, col_reg}<19'b0001011010111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0001011010111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0001011010111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0001011010111010000) && ({row_reg, col_reg}<19'b0001011010111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001011010111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0001011010111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0001011010111101010) && ({row_reg, col_reg}<19'b0001011100100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0001011100100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0001011100100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0001011100100111010) && ({row_reg, col_reg}<19'b0001011100100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001011100100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0001011100100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001011100100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0001011100100111111) && ({row_reg, col_reg}<19'b0001011100101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001011100101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0001011100101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0001011100101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0001011100101010100) && ({row_reg, col_reg}<19'b0001011100111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0001011100111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0001011100111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0001011100111010000) && ({row_reg, col_reg}<19'b0001011100111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001011100111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0001011100111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0001011100111101010) && ({row_reg, col_reg}<19'b0001011110100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0001011110100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0001011110100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0001011110100111010) && ({row_reg, col_reg}<19'b0001011110100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001011110100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0001011110100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001011110100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0001011110100111111) && ({row_reg, col_reg}<19'b0001011110101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001011110101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0001011110101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0001011110101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0001011110101010100) && ({row_reg, col_reg}<19'b0001011110111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0001011110111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0001011110111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0001011110111010000) && ({row_reg, col_reg}<19'b0001011110111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001011110111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0001011110111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0001011110111101010) && ({row_reg, col_reg}<19'b0001100000100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0001100000100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0001100000100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0001100000100111010) && ({row_reg, col_reg}<19'b0001100000100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001100000100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0001100000100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001100000100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0001100000100111111) && ({row_reg, col_reg}<19'b0001100000101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001100000101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0001100000101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0001100000101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0001100000101010100) && ({row_reg, col_reg}<19'b0001100000111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0001100000111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0001100000111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0001100000111010000) && ({row_reg, col_reg}<19'b0001100000111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001100000111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0001100000111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0001100000111101010) && ({row_reg, col_reg}<19'b0001100010100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0001100010100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0001100010100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0001100010100111010) && ({row_reg, col_reg}<19'b0001100010100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001100010100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0001100010100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001100010100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0001100010100111111) && ({row_reg, col_reg}<19'b0001100010101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001100010101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0001100010101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0001100010101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0001100010101010100) && ({row_reg, col_reg}<19'b0001100010111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0001100010111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0001100010111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0001100010111010000) && ({row_reg, col_reg}<19'b0001100010111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001100010111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0001100010111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0001100010111101010) && ({row_reg, col_reg}<19'b0001100100100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0001100100100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0001100100100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0001100100100111010) && ({row_reg, col_reg}<19'b0001100100100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001100100100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0001100100100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001100100100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0001100100100111111) && ({row_reg, col_reg}<19'b0001100100101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001100100101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0001100100101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0001100100101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0001100100101010100) && ({row_reg, col_reg}<19'b0001100100111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0001100100111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0001100100111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0001100100111010000) && ({row_reg, col_reg}<19'b0001100100111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001100100111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0001100100111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0001100100111101010) && ({row_reg, col_reg}<19'b0001100110100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0001100110100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0001100110100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0001100110100111010) && ({row_reg, col_reg}<19'b0001100110100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001100110100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0001100110100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001100110100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0001100110100111111) && ({row_reg, col_reg}<19'b0001100110101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001100110101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0001100110101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0001100110101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0001100110101010100) && ({row_reg, col_reg}<19'b0001100110111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0001100110111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0001100110111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0001100110111010000) && ({row_reg, col_reg}<19'b0001100110111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001100110111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0001100110111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0001100110111101010) && ({row_reg, col_reg}<19'b0001101000100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0001101000100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0001101000100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0001101000100111010) && ({row_reg, col_reg}<19'b0001101000100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001101000100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0001101000100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001101000100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0001101000100111111) && ({row_reg, col_reg}<19'b0001101000101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001101000101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0001101000101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0001101000101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0001101000101010100) && ({row_reg, col_reg}<19'b0001101000111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0001101000111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0001101000111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0001101000111010000) && ({row_reg, col_reg}<19'b0001101000111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001101000111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0001101000111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0001101000111101010) && ({row_reg, col_reg}<19'b0001101010100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0001101010100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0001101010100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0001101010100111010) && ({row_reg, col_reg}<19'b0001101010100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001101010100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0001101010100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001101010100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0001101010100111111) && ({row_reg, col_reg}<19'b0001101010101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001101010101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0001101010101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0001101010101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0001101010101010100) && ({row_reg, col_reg}<19'b0001101010111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0001101010111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0001101010111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0001101010111010000) && ({row_reg, col_reg}<19'b0001101010111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001101010111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0001101010111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0001101010111101010) && ({row_reg, col_reg}<19'b0001101100100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0001101100100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0001101100100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0001101100100111010) && ({row_reg, col_reg}<19'b0001101100100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001101100100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0001101100100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001101100100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0001101100100111111) && ({row_reg, col_reg}<19'b0001101100101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001101100101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0001101100101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0001101100101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0001101100101010100) && ({row_reg, col_reg}<19'b0001101100111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0001101100111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0001101100111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0001101100111010000) && ({row_reg, col_reg}<19'b0001101100111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001101100111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0001101100111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0001101100111101010) && ({row_reg, col_reg}<19'b0001101110100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0001101110100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0001101110100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0001101110100111010) && ({row_reg, col_reg}<19'b0001101110100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001101110100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0001101110100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001101110100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0001101110100111111) && ({row_reg, col_reg}<19'b0001101110101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001101110101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0001101110101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0001101110101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0001101110101010100) && ({row_reg, col_reg}<19'b0001101110111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0001101110111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0001101110111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0001101110111010000) && ({row_reg, col_reg}<19'b0001101110111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001101110111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0001101110111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0001101110111101010) && ({row_reg, col_reg}<19'b0001110000100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0001110000100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0001110000100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0001110000100111010) && ({row_reg, col_reg}<19'b0001110000100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001110000100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0001110000100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001110000100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0001110000100111111) && ({row_reg, col_reg}<19'b0001110000101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001110000101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0001110000101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0001110000101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0001110000101010100) && ({row_reg, col_reg}<19'b0001110000111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0001110000111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0001110000111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0001110000111010000) && ({row_reg, col_reg}<19'b0001110000111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001110000111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0001110000111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0001110000111101010) && ({row_reg, col_reg}<19'b0001110010100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0001110010100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0001110010100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0001110010100111010) && ({row_reg, col_reg}<19'b0001110010100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001110010100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0001110010100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001110010100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0001110010100111111) && ({row_reg, col_reg}<19'b0001110010101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001110010101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0001110010101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0001110010101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0001110010101010100) && ({row_reg, col_reg}<19'b0001110010111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0001110010111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0001110010111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0001110010111010000) && ({row_reg, col_reg}<19'b0001110010111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001110010111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0001110010111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0001110010111101010) && ({row_reg, col_reg}<19'b0001110100100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0001110100100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0001110100100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0001110100100111010) && ({row_reg, col_reg}<19'b0001110100100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001110100100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0001110100100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001110100100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0001110100100111111) && ({row_reg, col_reg}<19'b0001110100101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001110100101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0001110100101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0001110100101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0001110100101010100) && ({row_reg, col_reg}<19'b0001110100111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0001110100111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0001110100111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0001110100111010000) && ({row_reg, col_reg}<19'b0001110100111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001110100111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0001110100111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0001110100111101010) && ({row_reg, col_reg}<19'b0001110110100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0001110110100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0001110110100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0001110110100111010) && ({row_reg, col_reg}<19'b0001110110100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001110110100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0001110110100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001110110100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0001110110100111111) && ({row_reg, col_reg}<19'b0001110110101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001110110101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0001110110101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0001110110101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0001110110101010100) && ({row_reg, col_reg}<19'b0001110110111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0001110110111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0001110110111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0001110110111010000) && ({row_reg, col_reg}<19'b0001110110111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001110110111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0001110110111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0001110110111101010) && ({row_reg, col_reg}<19'b0001111000100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0001111000100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0001111000100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0001111000100111010) && ({row_reg, col_reg}<19'b0001111000100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001111000100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0001111000100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001111000100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0001111000100111111) && ({row_reg, col_reg}<19'b0001111000101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001111000101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0001111000101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0001111000101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0001111000101010100) && ({row_reg, col_reg}<19'b0001111000111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0001111000111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0001111000111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0001111000111010000) && ({row_reg, col_reg}<19'b0001111000111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001111000111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0001111000111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0001111000111101010) && ({row_reg, col_reg}<19'b0001111010100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0001111010100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0001111010100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0001111010100111010) && ({row_reg, col_reg}<19'b0001111010100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001111010100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0001111010100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001111010100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0001111010100111111) && ({row_reg, col_reg}<19'b0001111010101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001111010101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0001111010101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0001111010101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0001111010101010100) && ({row_reg, col_reg}<19'b0001111010111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0001111010111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0001111010111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0001111010111010000) && ({row_reg, col_reg}<19'b0001111010111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001111010111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0001111010111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0001111010111101010) && ({row_reg, col_reg}<19'b0001111100100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0001111100100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0001111100100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0001111100100111010) && ({row_reg, col_reg}<19'b0001111100100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001111100100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0001111100100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001111100100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0001111100100111111) && ({row_reg, col_reg}<19'b0001111100101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001111100101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0001111100101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0001111100101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0001111100101010100) && ({row_reg, col_reg}<19'b0001111100111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0001111100111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0001111100111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0001111100111010000) && ({row_reg, col_reg}<19'b0001111100111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001111100111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0001111100111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0001111100111101010) && ({row_reg, col_reg}<19'b0001111110100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0001111110100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0001111110100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0001111110100111010) && ({row_reg, col_reg}<19'b0001111110100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001111110100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0001111110100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001111110100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0001111110100111111) && ({row_reg, col_reg}<19'b0001111110101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001111110101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0001111110101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0001111110101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0001111110101010100) && ({row_reg, col_reg}<19'b0001111110111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0001111110111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0001111110111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0001111110111010000) && ({row_reg, col_reg}<19'b0001111110111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0001111110111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0001111110111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0001111110111101010) && ({row_reg, col_reg}<19'b0010000000100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010000000100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0010000000100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010000000100111010) && ({row_reg, col_reg}<19'b0010000000100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010000000100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0010000000100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010000000100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010000000100111111) && ({row_reg, col_reg}<19'b0010000000101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010000000101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0010000000101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0010000000101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0010000000101010100) && ({row_reg, col_reg}<19'b0010000000111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010000000111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0010000000111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010000000111010000) && ({row_reg, col_reg}<19'b0010000000111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010000000111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0010000000111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0010000000111101010) && ({row_reg, col_reg}<19'b0010000010100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010000010100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0010000010100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010000010100111010) && ({row_reg, col_reg}<19'b0010000010100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010000010100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0010000010100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010000010100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010000010100111111) && ({row_reg, col_reg}<19'b0010000010101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010000010101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0010000010101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0010000010101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0010000010101010100) && ({row_reg, col_reg}<19'b0010000010111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010000010111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0010000010111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010000010111010000) && ({row_reg, col_reg}<19'b0010000010111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010000010111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0010000010111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0010000010111101010) && ({row_reg, col_reg}<19'b0010000100100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010000100100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0010000100100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010000100100111010) && ({row_reg, col_reg}<19'b0010000100100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010000100100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0010000100100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010000100100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010000100100111111) && ({row_reg, col_reg}<19'b0010000100101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010000100101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0010000100101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0010000100101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0010000100101010100) && ({row_reg, col_reg}<19'b0010000100111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010000100111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0010000100111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010000100111010000) && ({row_reg, col_reg}<19'b0010000100111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010000100111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0010000100111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0010000100111101010) && ({row_reg, col_reg}<19'b0010000110100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010000110100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0010000110100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010000110100111010) && ({row_reg, col_reg}<19'b0010000110100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010000110100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0010000110100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010000110100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010000110100111111) && ({row_reg, col_reg}<19'b0010000110101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010000110101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0010000110101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0010000110101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0010000110101010100) && ({row_reg, col_reg}<19'b0010000110111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010000110111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0010000110111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010000110111010000) && ({row_reg, col_reg}<19'b0010000110111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010000110111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0010000110111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0010000110111101010) && ({row_reg, col_reg}<19'b0010001000100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010001000100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0010001000100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010001000100111010) && ({row_reg, col_reg}<19'b0010001000100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010001000100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0010001000100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010001000100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010001000100111111) && ({row_reg, col_reg}<19'b0010001000101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010001000101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0010001000101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0010001000101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0010001000101010100) && ({row_reg, col_reg}<19'b0010001000111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010001000111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0010001000111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010001000111010000) && ({row_reg, col_reg}<19'b0010001000111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010001000111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0010001000111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0010001000111101010) && ({row_reg, col_reg}<19'b0010001010100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010001010100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0010001010100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010001010100111010) && ({row_reg, col_reg}<19'b0010001010100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010001010100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0010001010100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010001010100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010001010100111111) && ({row_reg, col_reg}<19'b0010001010101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010001010101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0010001010101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0010001010101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0010001010101010100) && ({row_reg, col_reg}<19'b0010001010111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010001010111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0010001010111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010001010111010000) && ({row_reg, col_reg}<19'b0010001010111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010001010111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0010001010111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0010001010111101010) && ({row_reg, col_reg}<19'b0010001100100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010001100100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0010001100100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010001100100111010) && ({row_reg, col_reg}<19'b0010001100100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010001100100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0010001100100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010001100100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010001100100111111) && ({row_reg, col_reg}<19'b0010001100101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010001100101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0010001100101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0010001100101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0010001100101010100) && ({row_reg, col_reg}<19'b0010001100111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010001100111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0010001100111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010001100111010000) && ({row_reg, col_reg}<19'b0010001100111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010001100111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0010001100111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0010001100111101010) && ({row_reg, col_reg}<19'b0010001110100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010001110100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0010001110100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010001110100111010) && ({row_reg, col_reg}<19'b0010001110100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010001110100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0010001110100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010001110100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010001110100111111) && ({row_reg, col_reg}<19'b0010001110101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010001110101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0010001110101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0010001110101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0010001110101010100) && ({row_reg, col_reg}<19'b0010001110111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010001110111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0010001110111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010001110111010000) && ({row_reg, col_reg}<19'b0010001110111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010001110111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0010001110111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0010001110111101010) && ({row_reg, col_reg}<19'b0010010000100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010010000100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0010010000100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010010000100111010) && ({row_reg, col_reg}<19'b0010010000100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010010000100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0010010000100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010010000100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010010000100111111) && ({row_reg, col_reg}<19'b0010010000101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010010000101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0010010000101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0010010000101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0010010000101010100) && ({row_reg, col_reg}<19'b0010010000111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010010000111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0010010000111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010010000111010000) && ({row_reg, col_reg}<19'b0010010000111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010010000111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0010010000111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0010010000111101010) && ({row_reg, col_reg}<19'b0010010010100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010010010100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0010010010100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010010010100111010) && ({row_reg, col_reg}<19'b0010010010100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010010010100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0010010010100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010010010100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010010010100111111) && ({row_reg, col_reg}<19'b0010010010101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010010010101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0010010010101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0010010010101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0010010010101010100) && ({row_reg, col_reg}<19'b0010010010111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010010010111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0010010010111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010010010111010000) && ({row_reg, col_reg}<19'b0010010010111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010010010111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0010010010111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0010010010111101010) && ({row_reg, col_reg}<19'b0010010100100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010010100100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0010010100100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010010100100111010) && ({row_reg, col_reg}<19'b0010010100100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010010100100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0010010100100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010010100100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010010100100111111) && ({row_reg, col_reg}<19'b0010010100101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010010100101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0010010100101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0010010100101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0010010100101010100) && ({row_reg, col_reg}<19'b0010010100111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010010100111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0010010100111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010010100111010000) && ({row_reg, col_reg}<19'b0010010100111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010010100111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0010010100111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0010010100111101010) && ({row_reg, col_reg}<19'b0010010110100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010010110100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0010010110100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010010110100111010) && ({row_reg, col_reg}<19'b0010010110100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010010110100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0010010110100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010010110100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010010110100111111) && ({row_reg, col_reg}<19'b0010010110101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010010110101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0010010110101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0010010110101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0010010110101010100) && ({row_reg, col_reg}<19'b0010010110111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010010110111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0010010110111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010010110111010000) && ({row_reg, col_reg}<19'b0010010110111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010010110111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0010010110111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0010010110111101010) && ({row_reg, col_reg}<19'b0010011000100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010011000100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0010011000100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010011000100111010) && ({row_reg, col_reg}<19'b0010011000100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010011000100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0010011000100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010011000100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010011000100111111) && ({row_reg, col_reg}<19'b0010011000101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010011000101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0010011000101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0010011000101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0010011000101010100) && ({row_reg, col_reg}<19'b0010011000111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010011000111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0010011000111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010011000111010000) && ({row_reg, col_reg}<19'b0010011000111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010011000111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0010011000111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0010011000111101010) && ({row_reg, col_reg}<19'b0010011010100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010011010100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0010011010100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010011010100111010) && ({row_reg, col_reg}<19'b0010011010100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010011010100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0010011010100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010011010100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010011010100111111) && ({row_reg, col_reg}<19'b0010011010101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010011010101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0010011010101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0010011010101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0010011010101010100) && ({row_reg, col_reg}<19'b0010011010111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010011010111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0010011010111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010011010111010000) && ({row_reg, col_reg}<19'b0010011010111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010011010111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0010011010111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0010011010111101010) && ({row_reg, col_reg}<19'b0010011100100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010011100100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0010011100100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010011100100111010) && ({row_reg, col_reg}<19'b0010011100100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010011100100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0010011100100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010011100100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010011100100111111) && ({row_reg, col_reg}<19'b0010011100101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010011100101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0010011100101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0010011100101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0010011100101010100) && ({row_reg, col_reg}<19'b0010011100111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010011100111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0010011100111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010011100111010000) && ({row_reg, col_reg}<19'b0010011100111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010011100111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0010011100111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0010011100111101010) && ({row_reg, col_reg}<19'b0010011110100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010011110100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0010011110100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010011110100111010) && ({row_reg, col_reg}<19'b0010011110100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010011110100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0010011110100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010011110100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010011110100111111) && ({row_reg, col_reg}<19'b0010011110101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010011110101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0010011110101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0010011110101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0010011110101010100) && ({row_reg, col_reg}<19'b0010011110111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010011110111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0010011110111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010011110111010000) && ({row_reg, col_reg}<19'b0010011110111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010011110111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0010011110111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0010011110111101010) && ({row_reg, col_reg}<19'b0010100000100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010100000100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0010100000100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010100000100111010) && ({row_reg, col_reg}<19'b0010100000100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010100000100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0010100000100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010100000100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010100000100111111) && ({row_reg, col_reg}<19'b0010100000101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010100000101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0010100000101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0010100000101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0010100000101010100) && ({row_reg, col_reg}<19'b0010100000111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010100000111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0010100000111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010100000111010000) && ({row_reg, col_reg}<19'b0010100000111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010100000111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0010100000111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0010100000111101010) && ({row_reg, col_reg}<19'b0010100010100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010100010100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0010100010100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010100010100111010) && ({row_reg, col_reg}<19'b0010100010100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010100010100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0010100010100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010100010100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010100010100111111) && ({row_reg, col_reg}<19'b0010100010101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010100010101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0010100010101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0010100010101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0010100010101010100) && ({row_reg, col_reg}<19'b0010100010111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010100010111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0010100010111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010100010111010000) && ({row_reg, col_reg}<19'b0010100010111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010100010111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0010100010111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0010100010111101010) && ({row_reg, col_reg}<19'b0010100100100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010100100100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0010100100100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010100100100111010) && ({row_reg, col_reg}<19'b0010100100100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010100100100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0010100100100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010100100100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010100100100111111) && ({row_reg, col_reg}<19'b0010100100101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010100100101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0010100100101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0010100100101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0010100100101010100) && ({row_reg, col_reg}<19'b0010100100111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010100100111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0010100100111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010100100111010000) && ({row_reg, col_reg}<19'b0010100100111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010100100111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0010100100111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0010100100111101010) && ({row_reg, col_reg}<19'b0010100110100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010100110100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0010100110100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010100110100111010) && ({row_reg, col_reg}<19'b0010100110100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010100110100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0010100110100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010100110100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010100110100111111) && ({row_reg, col_reg}<19'b0010100110101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010100110101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0010100110101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0010100110101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0010100110101010100) && ({row_reg, col_reg}<19'b0010100110111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010100110111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0010100110111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010100110111010000) && ({row_reg, col_reg}<19'b0010100110111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010100110111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0010100110111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0010100110111101010) && ({row_reg, col_reg}<19'b0010101000100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010101000100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0010101000100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010101000100111010) && ({row_reg, col_reg}<19'b0010101000100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010101000100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0010101000100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010101000100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010101000100111111) && ({row_reg, col_reg}<19'b0010101000101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010101000101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0010101000101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0010101000101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0010101000101010100) && ({row_reg, col_reg}<19'b0010101000111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010101000111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0010101000111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010101000111010000) && ({row_reg, col_reg}<19'b0010101000111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010101000111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0010101000111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0010101000111101010) && ({row_reg, col_reg}<19'b0010101010100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010101010100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0010101010100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010101010100111010) && ({row_reg, col_reg}<19'b0010101010100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010101010100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0010101010100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010101010100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010101010100111111) && ({row_reg, col_reg}<19'b0010101010101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010101010101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0010101010101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0010101010101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0010101010101010100) && ({row_reg, col_reg}<19'b0010101010111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010101010111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0010101010111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010101010111010000) && ({row_reg, col_reg}<19'b0010101010111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010101010111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0010101010111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0010101010111101010) && ({row_reg, col_reg}<19'b0010101100100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010101100100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0010101100100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010101100100111010) && ({row_reg, col_reg}<19'b0010101100100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010101100100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0010101100100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010101100100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010101100100111111) && ({row_reg, col_reg}<19'b0010101100101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010101100101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0010101100101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0010101100101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0010101100101010100) && ({row_reg, col_reg}<19'b0010101100111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010101100111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0010101100111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010101100111010000) && ({row_reg, col_reg}<19'b0010101100111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010101100111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0010101100111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0010101100111101010) && ({row_reg, col_reg}<19'b0010101110100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010101110100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0010101110100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010101110100111010) && ({row_reg, col_reg}<19'b0010101110100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010101110100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0010101110100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010101110100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010101110100111111) && ({row_reg, col_reg}<19'b0010101110101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010101110101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0010101110101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0010101110101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0010101110101010100) && ({row_reg, col_reg}<19'b0010101110111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010101110111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0010101110111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010101110111010000) && ({row_reg, col_reg}<19'b0010101110111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010101110111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0010101110111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0010101110111101010) && ({row_reg, col_reg}<19'b0010110000100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010110000100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0010110000100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010110000100111010) && ({row_reg, col_reg}<19'b0010110000100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010110000100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0010110000100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010110000100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010110000100111111) && ({row_reg, col_reg}<19'b0010110000101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010110000101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0010110000101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0010110000101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0010110000101010100) && ({row_reg, col_reg}<19'b0010110000111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010110000111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0010110000111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010110000111010000) && ({row_reg, col_reg}<19'b0010110000111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010110000111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0010110000111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0010110000111101010) && ({row_reg, col_reg}<19'b0010110010100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010110010100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0010110010100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010110010100111010) && ({row_reg, col_reg}<19'b0010110010100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010110010100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0010110010100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010110010100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010110010100111111) && ({row_reg, col_reg}<19'b0010110010101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010110010101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0010110010101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0010110010101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0010110010101010100) && ({row_reg, col_reg}<19'b0010110010111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010110010111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0010110010111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010110010111010000) && ({row_reg, col_reg}<19'b0010110010111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010110010111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0010110010111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0010110010111101010) && ({row_reg, col_reg}<19'b0010110100100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010110100100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0010110100100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010110100100111010) && ({row_reg, col_reg}<19'b0010110100100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010110100100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0010110100100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010110100100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010110100100111111) && ({row_reg, col_reg}<19'b0010110100101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010110100101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0010110100101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0010110100101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0010110100101010100) && ({row_reg, col_reg}<19'b0010110100111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010110100111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0010110100111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010110100111010000) && ({row_reg, col_reg}<19'b0010110100111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010110100111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0010110100111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0010110100111101010) && ({row_reg, col_reg}<19'b0010110110100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010110110100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0010110110100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010110110100111010) && ({row_reg, col_reg}<19'b0010110110100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010110110100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0010110110100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010110110100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010110110100111111) && ({row_reg, col_reg}<19'b0010110110101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010110110101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0010110110101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0010110110101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0010110110101010100) && ({row_reg, col_reg}<19'b0010110110111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010110110111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0010110110111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010110110111010000) && ({row_reg, col_reg}<19'b0010110110111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010110110111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0010110110111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0010110110111101010) && ({row_reg, col_reg}<19'b0010111000100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010111000100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0010111000100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010111000100111010) && ({row_reg, col_reg}<19'b0010111000100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010111000100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0010111000100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010111000100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010111000100111111) && ({row_reg, col_reg}<19'b0010111000101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010111000101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0010111000101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0010111000101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0010111000101010100) && ({row_reg, col_reg}<19'b0010111000111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010111000111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0010111000111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010111000111010000) && ({row_reg, col_reg}<19'b0010111000111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010111000111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0010111000111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0010111000111101010) && ({row_reg, col_reg}<19'b0010111010100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010111010100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0010111010100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010111010100111010) && ({row_reg, col_reg}<19'b0010111010100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010111010100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0010111010100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010111010100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010111010100111111) && ({row_reg, col_reg}<19'b0010111010101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010111010101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0010111010101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0010111010101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0010111010101010100) && ({row_reg, col_reg}<19'b0010111010111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010111010111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0010111010111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010111010111010000) && ({row_reg, col_reg}<19'b0010111010111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010111010111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0010111010111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0010111010111101010) && ({row_reg, col_reg}<19'b0010111100100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010111100100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0010111100100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010111100100111010) && ({row_reg, col_reg}<19'b0010111100100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010111100100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0010111100100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010111100100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010111100100111111) && ({row_reg, col_reg}<19'b0010111100101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010111100101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0010111100101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0010111100101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0010111100101010100) && ({row_reg, col_reg}<19'b0010111100111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010111100111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0010111100111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010111100111010000) && ({row_reg, col_reg}<19'b0010111100111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010111100111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0010111100111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0010111100111101010) && ({row_reg, col_reg}<19'b0010111110100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010111110100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0010111110100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010111110100111010) && ({row_reg, col_reg}<19'b0010111110100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010111110100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0010111110100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010111110100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010111110100111111) && ({row_reg, col_reg}<19'b0010111110101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010111110101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0010111110101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0010111110101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0010111110101010100) && ({row_reg, col_reg}<19'b0010111110111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0010111110111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0010111110111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0010111110111010000) && ({row_reg, col_reg}<19'b0010111110111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0010111110111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0010111110111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0010111110111101010) && ({row_reg, col_reg}<19'b0011000000100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011000000100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0011000000100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011000000100111010) && ({row_reg, col_reg}<19'b0011000000100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011000000100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011000000100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011000000100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011000000100111111) && ({row_reg, col_reg}<19'b0011000000101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011000000101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011000000101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0011000000101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0011000000101010100) && ({row_reg, col_reg}<19'b0011000000111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011000000111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0011000000111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011000000111010000) && ({row_reg, col_reg}<19'b0011000000111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011000000111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0011000000111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0011000000111101010) && ({row_reg, col_reg}<19'b0011000010100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011000010100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0011000010100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011000010100111010) && ({row_reg, col_reg}<19'b0011000010100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011000010100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011000010100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011000010100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011000010100111111) && ({row_reg, col_reg}<19'b0011000010101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011000010101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011000010101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0011000010101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0011000010101010100) && ({row_reg, col_reg}<19'b0011000010111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011000010111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0011000010111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011000010111010000) && ({row_reg, col_reg}<19'b0011000010111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011000010111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0011000010111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0011000010111101010) && ({row_reg, col_reg}<19'b0011000100100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011000100100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0011000100100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011000100100111010) && ({row_reg, col_reg}<19'b0011000100100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011000100100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011000100100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011000100100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011000100100111111) && ({row_reg, col_reg}<19'b0011000100101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011000100101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011000100101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0011000100101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0011000100101010100) && ({row_reg, col_reg}<19'b0011000100111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011000100111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0011000100111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011000100111010000) && ({row_reg, col_reg}<19'b0011000100111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011000100111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0011000100111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0011000100111101010) && ({row_reg, col_reg}<19'b0011000110100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011000110100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0011000110100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011000110100111010) && ({row_reg, col_reg}<19'b0011000110100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011000110100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011000110100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011000110100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011000110100111111) && ({row_reg, col_reg}<19'b0011000110101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011000110101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011000110101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0011000110101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0011000110101010100) && ({row_reg, col_reg}<19'b0011000110111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011000110111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0011000110111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011000110111010000) && ({row_reg, col_reg}<19'b0011000110111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011000110111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0011000110111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0011000110111101010) && ({row_reg, col_reg}<19'b0011001000100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011001000100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0011001000100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011001000100111010) && ({row_reg, col_reg}<19'b0011001000100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011001000100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011001000100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011001000100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011001000100111111) && ({row_reg, col_reg}<19'b0011001000101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011001000101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011001000101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0011001000101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0011001000101010100) && ({row_reg, col_reg}<19'b0011001000111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011001000111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0011001000111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011001000111010000) && ({row_reg, col_reg}<19'b0011001000111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011001000111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0011001000111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0011001000111101010) && ({row_reg, col_reg}<19'b0011001010100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011001010100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0011001010100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011001010100111010) && ({row_reg, col_reg}<19'b0011001010100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011001010100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011001010100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011001010100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011001010100111111) && ({row_reg, col_reg}<19'b0011001010101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011001010101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011001010101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0011001010101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0011001010101010100) && ({row_reg, col_reg}<19'b0011001010111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011001010111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0011001010111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011001010111010000) && ({row_reg, col_reg}<19'b0011001010111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011001010111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0011001010111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0011001010111101010) && ({row_reg, col_reg}<19'b0011001100100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011001100100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0011001100100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011001100100111010) && ({row_reg, col_reg}<19'b0011001100100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011001100100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011001100100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011001100100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011001100100111111) && ({row_reg, col_reg}<19'b0011001100101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011001100101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011001100101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0011001100101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0011001100101010100) && ({row_reg, col_reg}<19'b0011001100111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011001100111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0011001100111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011001100111010000) && ({row_reg, col_reg}<19'b0011001100111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011001100111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0011001100111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0011001100111101010) && ({row_reg, col_reg}<19'b0011001110100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011001110100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0011001110100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011001110100111010) && ({row_reg, col_reg}<19'b0011001110100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011001110100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011001110100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011001110100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011001110100111111) && ({row_reg, col_reg}<19'b0011001110101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011001110101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011001110101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0011001110101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0011001110101010100) && ({row_reg, col_reg}<19'b0011001110111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011001110111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0011001110111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011001110111010000) && ({row_reg, col_reg}<19'b0011001110111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011001110111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0011001110111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0011001110111101010) && ({row_reg, col_reg}<19'b0011010000100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011010000100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0011010000100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011010000100111010) && ({row_reg, col_reg}<19'b0011010000100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011010000100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011010000100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011010000100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011010000100111111) && ({row_reg, col_reg}<19'b0011010000101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011010000101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011010000101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0011010000101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0011010000101010100) && ({row_reg, col_reg}<19'b0011010000111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011010000111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0011010000111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011010000111010000) && ({row_reg, col_reg}<19'b0011010000111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011010000111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0011010000111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0011010000111101010) && ({row_reg, col_reg}<19'b0011010010100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011010010100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0011010010100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011010010100111010) && ({row_reg, col_reg}<19'b0011010010100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011010010100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011010010100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011010010100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011010010100111111) && ({row_reg, col_reg}<19'b0011010010101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011010010101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011010010101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0011010010101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0011010010101010100) && ({row_reg, col_reg}<19'b0011010010111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011010010111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0011010010111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011010010111010000) && ({row_reg, col_reg}<19'b0011010010111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011010010111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0011010010111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0011010010111101010) && ({row_reg, col_reg}<19'b0011010100100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011010100100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0011010100100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011010100100111010) && ({row_reg, col_reg}<19'b0011010100100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011010100100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011010100100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011010100100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011010100100111111) && ({row_reg, col_reg}<19'b0011010100101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011010100101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011010100101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0011010100101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0011010100101010100) && ({row_reg, col_reg}<19'b0011010100111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011010100111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0011010100111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011010100111010000) && ({row_reg, col_reg}<19'b0011010100111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011010100111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0011010100111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0011010100111101010) && ({row_reg, col_reg}<19'b0011010110100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011010110100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0011010110100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011010110100111010) && ({row_reg, col_reg}<19'b0011010110100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011010110100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011010110100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011010110100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011010110100111111) && ({row_reg, col_reg}<19'b0011010110101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011010110101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011010110101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0011010110101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0011010110101010100) && ({row_reg, col_reg}<19'b0011010110111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011010110111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0011010110111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011010110111010000) && ({row_reg, col_reg}<19'b0011010110111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011010110111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0011010110111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0011010110111101010) && ({row_reg, col_reg}<19'b0011011000100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011011000100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0011011000100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011011000100111010) && ({row_reg, col_reg}<19'b0011011000100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011011000100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011011000100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011011000100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011011000100111111) && ({row_reg, col_reg}<19'b0011011000101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011011000101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011011000101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0011011000101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0011011000101010100) && ({row_reg, col_reg}<19'b0011011000111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011011000111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0011011000111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011011000111010000) && ({row_reg, col_reg}<19'b0011011000111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011011000111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0011011000111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0011011000111101010) && ({row_reg, col_reg}<19'b0011011010100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011011010100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0011011010100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011011010100111010) && ({row_reg, col_reg}<19'b0011011010100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011011010100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011011010100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011011010100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011011010100111111) && ({row_reg, col_reg}<19'b0011011010101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011011010101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011011010101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0011011010101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0011011010101010100) && ({row_reg, col_reg}<19'b0011011010111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011011010111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0011011010111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011011010111010000) && ({row_reg, col_reg}<19'b0011011010111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011011010111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0011011010111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0011011010111101010) && ({row_reg, col_reg}<19'b0011011100100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011011100100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0011011100100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011011100100111010) && ({row_reg, col_reg}<19'b0011011100100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011011100100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011011100100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011011100100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011011100100111111) && ({row_reg, col_reg}<19'b0011011100101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011011100101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011011100101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0011011100101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0011011100101010100) && ({row_reg, col_reg}<19'b0011011100111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011011100111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0011011100111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011011100111010000) && ({row_reg, col_reg}<19'b0011011100111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011011100111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0011011100111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0011011100111101010) && ({row_reg, col_reg}<19'b0011011110100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011011110100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0011011110100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011011110100111010) && ({row_reg, col_reg}<19'b0011011110100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011011110100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011011110100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011011110100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011011110100111111) && ({row_reg, col_reg}<19'b0011011110101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011011110101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011011110101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0011011110101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0011011110101010100) && ({row_reg, col_reg}<19'b0011011110111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011011110111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0011011110111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011011110111010000) && ({row_reg, col_reg}<19'b0011011110111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011011110111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0011011110111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0011011110111101010) && ({row_reg, col_reg}<19'b0011100000100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011100000100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0011100000100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011100000100111010) && ({row_reg, col_reg}<19'b0011100000100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011100000100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011100000100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011100000100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011100000100111111) && ({row_reg, col_reg}<19'b0011100000101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011100000101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011100000101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0011100000101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0011100000101010100) && ({row_reg, col_reg}<19'b0011100000111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011100000111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0011100000111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011100000111010000) && ({row_reg, col_reg}<19'b0011100000111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011100000111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0011100000111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0011100000111101010) && ({row_reg, col_reg}<19'b0011100010100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011100010100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0011100010100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011100010100111010) && ({row_reg, col_reg}<19'b0011100010100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011100010100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011100010100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011100010100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011100010100111111) && ({row_reg, col_reg}<19'b0011100010101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011100010101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011100010101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0011100010101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0011100010101010100) && ({row_reg, col_reg}<19'b0011100010111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011100010111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0011100010111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011100010111010000) && ({row_reg, col_reg}<19'b0011100010111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011100010111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0011100010111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0011100010111101010) && ({row_reg, col_reg}<19'b0011100100100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011100100100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0011100100100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011100100100111010) && ({row_reg, col_reg}<19'b0011100100100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011100100100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011100100100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011100100100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011100100100111111) && ({row_reg, col_reg}<19'b0011100100101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011100100101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011100100101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0011100100101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0011100100101010100) && ({row_reg, col_reg}<19'b0011100100111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011100100111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0011100100111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011100100111010000) && ({row_reg, col_reg}<19'b0011100100111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011100100111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0011100100111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0011100100111101010) && ({row_reg, col_reg}<19'b0011100110100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011100110100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0011100110100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011100110100111010) && ({row_reg, col_reg}<19'b0011100110100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011100110100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011100110100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011100110100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011100110100111111) && ({row_reg, col_reg}<19'b0011100110101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011100110101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011100110101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0011100110101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0011100110101010100) && ({row_reg, col_reg}<19'b0011100110111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011100110111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0011100110111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011100110111010000) && ({row_reg, col_reg}<19'b0011100110111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011100110111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0011100110111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0011100110111101010) && ({row_reg, col_reg}<19'b0011101000100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011101000100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0011101000100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011101000100111010) && ({row_reg, col_reg}<19'b0011101000100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011101000100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011101000100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011101000100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011101000100111111) && ({row_reg, col_reg}<19'b0011101000101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011101000101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011101000101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0011101000101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0011101000101010100) && ({row_reg, col_reg}<19'b0011101000111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011101000111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0011101000111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011101000111010000) && ({row_reg, col_reg}<19'b0011101000111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011101000111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0011101000111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0011101000111101010) && ({row_reg, col_reg}<19'b0011101010100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011101010100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0011101010100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011101010100111010) && ({row_reg, col_reg}<19'b0011101010100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011101010100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011101010100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011101010100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011101010100111111) && ({row_reg, col_reg}<19'b0011101010101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011101010101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011101010101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0011101010101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0011101010101010100) && ({row_reg, col_reg}<19'b0011101010111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011101010111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0011101010111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011101010111010000) && ({row_reg, col_reg}<19'b0011101010111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011101010111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0011101010111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0011101010111101010) && ({row_reg, col_reg}<19'b0011101100100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011101100100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0011101100100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011101100100111010) && ({row_reg, col_reg}<19'b0011101100100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011101100100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011101100100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011101100100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011101100100111111) && ({row_reg, col_reg}<19'b0011101100101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011101100101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011101100101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0011101100101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0011101100101010100) && ({row_reg, col_reg}<19'b0011101100111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011101100111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0011101100111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011101100111010000) && ({row_reg, col_reg}<19'b0011101100111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011101100111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0011101100111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0011101100111101010) && ({row_reg, col_reg}<19'b0011101110100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011101110100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0011101110100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011101110100111010) && ({row_reg, col_reg}<19'b0011101110100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011101110100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011101110100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011101110100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011101110100111111) && ({row_reg, col_reg}<19'b0011101110101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011101110101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011101110101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0011101110101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0011101110101010100) && ({row_reg, col_reg}<19'b0011101110111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011101110111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0011101110111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011101110111010000) && ({row_reg, col_reg}<19'b0011101110111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011101110111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0011101110111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0011101110111101010) && ({row_reg, col_reg}<19'b0011110000100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011110000100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0011110000100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011110000100111010) && ({row_reg, col_reg}<19'b0011110000100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011110000100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011110000100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011110000100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011110000100111111) && ({row_reg, col_reg}<19'b0011110000101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011110000101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011110000101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0011110000101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0011110000101010100) && ({row_reg, col_reg}<19'b0011110000111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011110000111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0011110000111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011110000111010000) && ({row_reg, col_reg}<19'b0011110000111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011110000111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0011110000111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0011110000111101010) && ({row_reg, col_reg}<19'b0011110010100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011110010100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0011110010100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011110010100111010) && ({row_reg, col_reg}<19'b0011110010100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011110010100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011110010100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011110010100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011110010100111111) && ({row_reg, col_reg}<19'b0011110010101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011110010101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011110010101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0011110010101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0011110010101010100) && ({row_reg, col_reg}<19'b0011110010111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011110010111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0011110010111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011110010111010000) && ({row_reg, col_reg}<19'b0011110010111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011110010111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0011110010111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0011110010111101010) && ({row_reg, col_reg}<19'b0011110100100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011110100100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0011110100100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011110100100111010) && ({row_reg, col_reg}<19'b0011110100100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011110100100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011110100100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011110100100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011110100100111111) && ({row_reg, col_reg}<19'b0011110100101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011110100101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011110100101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0011110100101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0011110100101010100) && ({row_reg, col_reg}<19'b0011110100111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011110100111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0011110100111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011110100111010000) && ({row_reg, col_reg}<19'b0011110100111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011110100111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0011110100111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0011110100111101010) && ({row_reg, col_reg}<19'b0011110110100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011110110100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0011110110100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011110110100111010) && ({row_reg, col_reg}<19'b0011110110100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011110110100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011110110100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011110110100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011110110100111111) && ({row_reg, col_reg}<19'b0011110110101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011110110101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011110110101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0011110110101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0011110110101010100) && ({row_reg, col_reg}<19'b0011110110111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011110110111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0011110110111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011110110111010000) && ({row_reg, col_reg}<19'b0011110110111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011110110111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0011110110111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0011110110111101010) && ({row_reg, col_reg}<19'b0011111000100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011111000100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0011111000100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011111000100111010) && ({row_reg, col_reg}<19'b0011111000100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011111000100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011111000100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011111000100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011111000100111111) && ({row_reg, col_reg}<19'b0011111000101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011111000101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011111000101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0011111000101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0011111000101010100) && ({row_reg, col_reg}<19'b0011111000111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011111000111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0011111000111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011111000111010000) && ({row_reg, col_reg}<19'b0011111000111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011111000111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0011111000111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0011111000111101010) && ({row_reg, col_reg}<19'b0011111010100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011111010100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0011111010100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011111010100111010) && ({row_reg, col_reg}<19'b0011111010100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011111010100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011111010100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011111010100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011111010100111111) && ({row_reg, col_reg}<19'b0011111010101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011111010101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011111010101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0011111010101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0011111010101010100) && ({row_reg, col_reg}<19'b0011111010111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011111010111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0011111010111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011111010111010000) && ({row_reg, col_reg}<19'b0011111010111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011111010111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0011111010111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0011111010111101010) && ({row_reg, col_reg}<19'b0011111100100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011111100100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0011111100100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011111100100111010) && ({row_reg, col_reg}<19'b0011111100100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011111100100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011111100100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011111100100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011111100100111111) && ({row_reg, col_reg}<19'b0011111100101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011111100101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011111100101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0011111100101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0011111100101010100) && ({row_reg, col_reg}<19'b0011111100111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011111100111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0011111100111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011111100111010000) && ({row_reg, col_reg}<19'b0011111100111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011111100111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0011111100111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0011111100111101010) && ({row_reg, col_reg}<19'b0011111110100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011111110100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0011111110100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011111110100111010) && ({row_reg, col_reg}<19'b0011111110100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011111110100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011111110100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011111110100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011111110100111111) && ({row_reg, col_reg}<19'b0011111110101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011111110101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0011111110101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0011111110101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0011111110101010100) && ({row_reg, col_reg}<19'b0011111110111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0011111110111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0011111110111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0011111110111010000) && ({row_reg, col_reg}<19'b0011111110111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0011111110111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0011111110111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0011111110111101010) && ({row_reg, col_reg}<19'b0100000000100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100000000100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0100000000100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100000000100111010) && ({row_reg, col_reg}<19'b0100000000100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100000000100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0100000000100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100000000100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100000000100111111) && ({row_reg, col_reg}<19'b0100000000101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100000000101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0100000000101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0100000000101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0100000000101010100) && ({row_reg, col_reg}<19'b0100000000111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100000000111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0100000000111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100000000111010000) && ({row_reg, col_reg}<19'b0100000000111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100000000111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0100000000111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0100000000111101010) && ({row_reg, col_reg}<19'b0100000010100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100000010100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0100000010100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100000010100111010) && ({row_reg, col_reg}<19'b0100000010100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100000010100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0100000010100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100000010100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100000010100111111) && ({row_reg, col_reg}<19'b0100000010101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100000010101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0100000010101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0100000010101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0100000010101010100) && ({row_reg, col_reg}<19'b0100000010111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100000010111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0100000010111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100000010111010000) && ({row_reg, col_reg}<19'b0100000010111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100000010111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0100000010111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0100000010111101010) && ({row_reg, col_reg}<19'b0100000100100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100000100100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0100000100100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100000100100111010) && ({row_reg, col_reg}<19'b0100000100100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100000100100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0100000100100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100000100100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100000100100111111) && ({row_reg, col_reg}<19'b0100000100101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100000100101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0100000100101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0100000100101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0100000100101010100) && ({row_reg, col_reg}<19'b0100000100111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100000100111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0100000100111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100000100111010000) && ({row_reg, col_reg}<19'b0100000100111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100000100111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0100000100111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0100000100111101010) && ({row_reg, col_reg}<19'b0100000110100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100000110100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0100000110100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100000110100111010) && ({row_reg, col_reg}<19'b0100000110100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100000110100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0100000110100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100000110100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100000110100111111) && ({row_reg, col_reg}<19'b0100000110101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100000110101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0100000110101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0100000110101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0100000110101010100) && ({row_reg, col_reg}<19'b0100000110111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100000110111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0100000110111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100000110111010000) && ({row_reg, col_reg}<19'b0100000110111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100000110111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0100000110111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0100000110111101010) && ({row_reg, col_reg}<19'b0100001000100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100001000100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0100001000100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100001000100111010) && ({row_reg, col_reg}<19'b0100001000100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100001000100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0100001000100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100001000100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100001000100111111) && ({row_reg, col_reg}<19'b0100001000101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100001000101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0100001000101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0100001000101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0100001000101010100) && ({row_reg, col_reg}<19'b0100001000111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100001000111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0100001000111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100001000111010000) && ({row_reg, col_reg}<19'b0100001000111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100001000111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0100001000111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0100001000111101010) && ({row_reg, col_reg}<19'b0100001010100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100001010100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0100001010100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100001010100111010) && ({row_reg, col_reg}<19'b0100001010100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100001010100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0100001010100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100001010100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100001010100111111) && ({row_reg, col_reg}<19'b0100001010101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100001010101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0100001010101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0100001010101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0100001010101010100) && ({row_reg, col_reg}<19'b0100001010111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100001010111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0100001010111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100001010111010000) && ({row_reg, col_reg}<19'b0100001010111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100001010111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0100001010111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0100001010111101010) && ({row_reg, col_reg}<19'b0100001100100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100001100100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0100001100100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100001100100111010) && ({row_reg, col_reg}<19'b0100001100100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100001100100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0100001100100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100001100100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100001100100111111) && ({row_reg, col_reg}<19'b0100001100101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100001100101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0100001100101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0100001100101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0100001100101010100) && ({row_reg, col_reg}<19'b0100001100111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100001100111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0100001100111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100001100111010000) && ({row_reg, col_reg}<19'b0100001100111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100001100111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0100001100111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0100001100111101010) && ({row_reg, col_reg}<19'b0100001110100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100001110100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0100001110100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100001110100111010) && ({row_reg, col_reg}<19'b0100001110100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100001110100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0100001110100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100001110100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100001110100111111) && ({row_reg, col_reg}<19'b0100001110101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100001110101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0100001110101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0100001110101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0100001110101010100) && ({row_reg, col_reg}<19'b0100001110111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100001110111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0100001110111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100001110111010000) && ({row_reg, col_reg}<19'b0100001110111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100001110111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0100001110111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0100001110111101010) && ({row_reg, col_reg}<19'b0100010000100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100010000100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0100010000100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100010000100111010) && ({row_reg, col_reg}<19'b0100010000100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100010000100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0100010000100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100010000100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100010000100111111) && ({row_reg, col_reg}<19'b0100010000101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100010000101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0100010000101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0100010000101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0100010000101010100) && ({row_reg, col_reg}<19'b0100010000111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100010000111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0100010000111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100010000111010000) && ({row_reg, col_reg}<19'b0100010000111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100010000111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0100010000111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0100010000111101010) && ({row_reg, col_reg}<19'b0100010010100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100010010100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0100010010100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100010010100111010) && ({row_reg, col_reg}<19'b0100010010100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100010010100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0100010010100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100010010100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100010010100111111) && ({row_reg, col_reg}<19'b0100010010101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100010010101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0100010010101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0100010010101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0100010010101010100) && ({row_reg, col_reg}<19'b0100010010111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100010010111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0100010010111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100010010111010000) && ({row_reg, col_reg}<19'b0100010010111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100010010111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0100010010111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0100010010111101010) && ({row_reg, col_reg}<19'b0100010100100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100010100100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0100010100100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100010100100111010) && ({row_reg, col_reg}<19'b0100010100100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100010100100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0100010100100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100010100100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100010100100111111) && ({row_reg, col_reg}<19'b0100010100101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100010100101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0100010100101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0100010100101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0100010100101010100) && ({row_reg, col_reg}<19'b0100010100111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100010100111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0100010100111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100010100111010000) && ({row_reg, col_reg}<19'b0100010100111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100010100111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0100010100111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0100010100111101010) && ({row_reg, col_reg}<19'b0100010110100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100010110100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0100010110100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100010110100111010) && ({row_reg, col_reg}<19'b0100010110100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100010110100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0100010110100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100010110100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100010110100111111) && ({row_reg, col_reg}<19'b0100010110101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100010110101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0100010110101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0100010110101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0100010110101010100) && ({row_reg, col_reg}<19'b0100010110111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100010110111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0100010110111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100010110111010000) && ({row_reg, col_reg}<19'b0100010110111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100010110111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0100010110111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0100010110111101010) && ({row_reg, col_reg}<19'b0100011000100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100011000100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0100011000100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100011000100111010) && ({row_reg, col_reg}<19'b0100011000100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100011000100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0100011000100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100011000100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100011000100111111) && ({row_reg, col_reg}<19'b0100011000101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100011000101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0100011000101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0100011000101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0100011000101010100) && ({row_reg, col_reg}<19'b0100011000111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100011000111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0100011000111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100011000111010000) && ({row_reg, col_reg}<19'b0100011000111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100011000111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0100011000111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0100011000111101010) && ({row_reg, col_reg}<19'b0100011010100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100011010100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0100011010100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100011010100111010) && ({row_reg, col_reg}<19'b0100011010100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100011010100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0100011010100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100011010100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100011010100111111) && ({row_reg, col_reg}<19'b0100011010101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100011010101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0100011010101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0100011010101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0100011010101010100) && ({row_reg, col_reg}<19'b0100011010111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100011010111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0100011010111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100011010111010000) && ({row_reg, col_reg}<19'b0100011010111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100011010111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0100011010111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0100011010111101010) && ({row_reg, col_reg}<19'b0100011100100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100011100100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0100011100100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100011100100111010) && ({row_reg, col_reg}<19'b0100011100100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100011100100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0100011100100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100011100100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100011100100111111) && ({row_reg, col_reg}<19'b0100011100101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100011100101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0100011100101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0100011100101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0100011100101010100) && ({row_reg, col_reg}<19'b0100011100111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100011100111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0100011100111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100011100111010000) && ({row_reg, col_reg}<19'b0100011100111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100011100111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0100011100111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0100011100111101010) && ({row_reg, col_reg}<19'b0100011110100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100011110100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0100011110100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100011110100111010) && ({row_reg, col_reg}<19'b0100011110100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100011110100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0100011110100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100011110100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100011110100111111) && ({row_reg, col_reg}<19'b0100011110101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100011110101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0100011110101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0100011110101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0100011110101010100) && ({row_reg, col_reg}<19'b0100011110111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100011110111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0100011110111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100011110111010000) && ({row_reg, col_reg}<19'b0100011110111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100011110111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0100011110111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0100011110111101010) && ({row_reg, col_reg}<19'b0100100000100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100100000100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0100100000100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100100000100111010) && ({row_reg, col_reg}<19'b0100100000100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100100000100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0100100000100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100100000100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100100000100111111) && ({row_reg, col_reg}<19'b0100100000101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100100000101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0100100000101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0100100000101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0100100000101010100) && ({row_reg, col_reg}<19'b0100100000111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100100000111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0100100000111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100100000111010000) && ({row_reg, col_reg}<19'b0100100000111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100100000111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0100100000111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0100100000111101010) && ({row_reg, col_reg}<19'b0100100010100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100100010100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0100100010100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100100010100111010) && ({row_reg, col_reg}<19'b0100100010100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100100010100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0100100010100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100100010100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100100010100111111) && ({row_reg, col_reg}<19'b0100100010101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100100010101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0100100010101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0100100010101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0100100010101010100) && ({row_reg, col_reg}<19'b0100100010111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100100010111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0100100010111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100100010111010000) && ({row_reg, col_reg}<19'b0100100010111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100100010111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0100100010111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0100100010111101010) && ({row_reg, col_reg}<19'b0100100100100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100100100100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0100100100100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100100100100111010) && ({row_reg, col_reg}<19'b0100100100100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100100100100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0100100100100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100100100100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100100100100111111) && ({row_reg, col_reg}<19'b0100100100101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100100100101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0100100100101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0100100100101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0100100100101010100) && ({row_reg, col_reg}<19'b0100100100111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100100100111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0100100100111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100100100111010000) && ({row_reg, col_reg}<19'b0100100100111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100100100111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0100100100111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0100100100111101010) && ({row_reg, col_reg}<19'b0100100110100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100100110100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0100100110100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100100110100111010) && ({row_reg, col_reg}<19'b0100100110100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100100110100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0100100110100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100100110100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100100110100111111) && ({row_reg, col_reg}<19'b0100100110101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100100110101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0100100110101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0100100110101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0100100110101010100) && ({row_reg, col_reg}<19'b0100100110111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100100110111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0100100110111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100100110111010000) && ({row_reg, col_reg}<19'b0100100110111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100100110111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0100100110111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0100100110111101010) && ({row_reg, col_reg}<19'b0100101000100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100101000100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0100101000100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100101000100111010) && ({row_reg, col_reg}<19'b0100101000100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100101000100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0100101000100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100101000100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100101000100111111) && ({row_reg, col_reg}<19'b0100101000101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100101000101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0100101000101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0100101000101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0100101000101010100) && ({row_reg, col_reg}<19'b0100101000111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100101000111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0100101000111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100101000111010000) && ({row_reg, col_reg}<19'b0100101000111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100101000111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0100101000111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0100101000111101010) && ({row_reg, col_reg}<19'b0100101010100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100101010100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0100101010100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100101010100111010) && ({row_reg, col_reg}<19'b0100101010100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100101010100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0100101010100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100101010100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100101010100111111) && ({row_reg, col_reg}<19'b0100101010101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100101010101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0100101010101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0100101010101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0100101010101010100) && ({row_reg, col_reg}<19'b0100101010111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100101010111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0100101010111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100101010111010000) && ({row_reg, col_reg}<19'b0100101010111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100101010111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0100101010111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0100101010111101010) && ({row_reg, col_reg}<19'b0100101100100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100101100100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0100101100100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100101100100111010) && ({row_reg, col_reg}<19'b0100101100100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100101100100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0100101100100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100101100100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100101100100111111) && ({row_reg, col_reg}<19'b0100101100101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100101100101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0100101100101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0100101100101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0100101100101010100) && ({row_reg, col_reg}<19'b0100101100111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100101100111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0100101100111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100101100111010000) && ({row_reg, col_reg}<19'b0100101100111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100101100111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0100101100111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0100101100111101010) && ({row_reg, col_reg}<19'b0100101110100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100101110100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0100101110100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100101110100111010) && ({row_reg, col_reg}<19'b0100101110100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100101110100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0100101110100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100101110100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100101110100111111) && ({row_reg, col_reg}<19'b0100101110101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100101110101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0100101110101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0100101110101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0100101110101010100) && ({row_reg, col_reg}<19'b0100101110111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100101110111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0100101110111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100101110111010000) && ({row_reg, col_reg}<19'b0100101110111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100101110111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0100101110111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0100101110111101010) && ({row_reg, col_reg}<19'b0100110000100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100110000100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0100110000100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100110000100111010) && ({row_reg, col_reg}<19'b0100110000100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100110000100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0100110000100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100110000100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100110000100111111) && ({row_reg, col_reg}<19'b0100110000101010000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0100110000101010000) && ({row_reg, col_reg}<19'b0100110000101010010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0100110000101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0100110000101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0100110000101010100) && ({row_reg, col_reg}<19'b0100110000111001101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100110000111001101)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0100110000111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0100110000111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100110000111010000) && ({row_reg, col_reg}<19'b0100110000111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100110000111101000)) color_data = 12'b101010101010;

		if(({row_reg, col_reg}>=19'b0100110000111101001) && ({row_reg, col_reg}<19'b0100110010100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100110010100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0100110010100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100110010100111010) && ({row_reg, col_reg}<19'b0100110010100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100110010100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0100110010100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100110010100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100110010100111111) && ({row_reg, col_reg}<19'b0100110010101010010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100110010101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0100110010101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0100110010101010100) && ({row_reg, col_reg}<19'b0100110010111001101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100110010111001101)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0100110010111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0100110010111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100110010111010000) && ({row_reg, col_reg}<19'b0100110010111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100110010111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0100110010111101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=19'b0100110010111101010) && ({row_reg, col_reg}<19'b0100110011001111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100110011001111000)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0100110011001111001) && ({row_reg, col_reg}<19'b0100110100010101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100110100010101100)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=19'b0100110100010101101) && ({row_reg, col_reg}<19'b0100110100010110000)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0100110100010110000) && ({row_reg, col_reg}<19'b0100110100100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0100110100100111000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0100110100100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100110100100111010) && ({row_reg, col_reg}<19'b0100110100100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100110100100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0100110100100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100110100100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100110100100111111) && ({row_reg, col_reg}<19'b0100110100101010000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0100110100101010000) && ({row_reg, col_reg}<19'b0100110100101010010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0100110100101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0100110100101010011)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=19'b0100110100101010100) && ({row_reg, col_reg}<19'b0100110100111001100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0100110100111001100)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0100110100111001101)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0100110100111001110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0100110100111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100110100111010000) && ({row_reg, col_reg}<19'b0100110100111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100110100111101000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=19'b0100110100111101001) && ({row_reg, col_reg}<19'b0100110101001110011)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=19'b0100110101001110011) && ({row_reg, col_reg}<19'b0100110101001110101)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0100110101001110101)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0100110101001110110) && ({row_reg, col_reg}<19'b0100110110010101001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100110110010101001)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0100110110010101010) && ({row_reg, col_reg}<19'b0100110110010101100)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0100110110010101100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=19'b0100110110010101101) && ({row_reg, col_reg}<19'b0100110110010101111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=19'b0100110110010101111) && ({row_reg, col_reg}<19'b0100110110100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0100110110100111001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100110110100111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0100110110100111011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100110110100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100110110100111101) && ({row_reg, col_reg}<19'b0100110110100111111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100110110100111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100110110101000000) && ({row_reg, col_reg}<19'b0100110110101010011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0100110110101010011) && ({row_reg, col_reg}<19'b0100110110111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100110110111001111) && ({row_reg, col_reg}<19'b0100110110111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100110110111101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0100110110111101001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=19'b0100110110111101010) && ({row_reg, col_reg}<19'b0100110110111101101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100110110111101101) && ({row_reg, col_reg}<19'b0100110110111101111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=19'b0100110110111101111) && ({row_reg, col_reg}<19'b0100110111001110011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100110111001110011) && ({row_reg, col_reg}<19'b0100110111001110101)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0100110111001110101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0100110111001110110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0100110111001110111)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0100110111001111000)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0100110111001111001) && ({row_reg, col_reg}<19'b0100111000010100111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100111000010100111)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0100111000010101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0100111000010101001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=19'b0100111000010101010) && ({row_reg, col_reg}<19'b0100111000010101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100111000010101100) && ({row_reg, col_reg}<19'b0100111000010101110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0100111000010101110) && ({row_reg, col_reg}<19'b0100111000010110000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100111000010110000) && ({row_reg, col_reg}<19'b0100111000100111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100111000100111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100111000100111011) && ({row_reg, col_reg}<19'b0100111000101010000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0100111000101010000) && ({row_reg, col_reg}<19'b0100111000101010010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0100111000101010010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100111000101010011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0100111000101010100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0100111000101010101) && ({row_reg, col_reg}<19'b0100111000101011000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100111000101011000) && ({row_reg, col_reg}<19'b0100111000111001000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0100111000111001000) && ({row_reg, col_reg}<19'b0100111000111001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0100111000111001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0100111000111001101) && ({row_reg, col_reg}<19'b0100111000111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100111000111001111) && ({row_reg, col_reg}<19'b0100111000111101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100111000111101101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100111000111101110) && ({row_reg, col_reg}<19'b0100111001001110000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100111001001110000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100111001001110001) && ({row_reg, col_reg}<19'b0100111001001110011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100111001001110011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100111001001110100) && ({row_reg, col_reg}<19'b0100111001001110110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0100111001001110110) && ({row_reg, col_reg}<19'b0100111001001111000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0100111001001111000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0100111001001111001)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=19'b0100111001001111010) && ({row_reg, col_reg}<19'b0100111010010100101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100111010010100101)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0100111010010100110)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0100111010010100111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0100111010010101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100111010010101001) && ({row_reg, col_reg}<19'b0100111010010101011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0100111010010101011) && ({row_reg, col_reg}<19'b0100111010010101111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100111010010101111) && ({row_reg, col_reg}<19'b0100111010100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0100111010100111101) && ({row_reg, col_reg}<19'b0100111010100111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100111010100111111) && ({row_reg, col_reg}<19'b0100111010101010000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0100111010101010000) && ({row_reg, col_reg}<19'b0100111010101010010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100111010101010010) && ({row_reg, col_reg}<19'b0100111010111001011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100111010111001011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0100111010111001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0100111010111001101) && ({row_reg, col_reg}<19'b0100111010111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100111010111001111) && ({row_reg, col_reg}<19'b0100111010111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0100111010111101000) && ({row_reg, col_reg}<19'b0100111010111101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100111010111101100) && ({row_reg, col_reg}<19'b0100111010111101111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100111010111101111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100111010111110000) && ({row_reg, col_reg}<19'b0100111011001110100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100111011001110100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100111011001110101) && ({row_reg, col_reg}<19'b0100111011001111001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100111011001111001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0100111011001111010)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0100111011001111011)) color_data = 12'b110111011101;

		if(({row_reg, col_reg}>=19'b0100111011001111100) && ({row_reg, col_reg}<19'b0100111100010100100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100111100010100100)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0100111100010100101)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0100111100010100110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=19'b0100111100010100111) && ({row_reg, col_reg}<19'b0100111100010101110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100111100010101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100111100010101111) && ({row_reg, col_reg}<19'b0100111100100111000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100111100100111000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100111100100111001) && ({row_reg, col_reg}<19'b0100111100100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0100111100100111101) && ({row_reg, col_reg}<19'b0100111100100111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100111100100111111) && ({row_reg, col_reg}<19'b0100111100101010010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100111100101010010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0100111100101010011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0100111100101010100) && ({row_reg, col_reg}<19'b0100111100101011000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100111100101011000) && ({row_reg, col_reg}<19'b0100111100111001000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0100111100111001000) && ({row_reg, col_reg}<19'b0100111100111001010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0100111100111001010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100111100111001011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100111100111001100) && ({row_reg, col_reg}<19'b0100111100111101010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100111100111101010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100111100111101011) && ({row_reg, col_reg}<19'b0100111100111101111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100111100111101111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100111100111110000) && ({row_reg, col_reg}<19'b0100111101001110000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0100111101001110000) && ({row_reg, col_reg}<19'b0100111101001110011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100111101001110011) && ({row_reg, col_reg}<19'b0100111101001111000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100111101001111000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0100111101001111001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100111101001111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0100111101001111011)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0100111101001111100)) color_data = 12'b110111011101;

		if(({row_reg, col_reg}>=19'b0100111101001111101) && ({row_reg, col_reg}<19'b0100111110010100100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0100111110010100100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0100111110010100101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0100111110010100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100111110010100111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0100111110010101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0100111110010101001) && ({row_reg, col_reg}<19'b0100111110010101101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100111110010101101) && ({row_reg, col_reg}<19'b0100111110100111001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100111110100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0100111110100111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100111110100111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100111110100111100) && ({row_reg, col_reg}<19'b0100111110101010000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100111110101010000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100111110101010001) && ({row_reg, col_reg}<19'b0100111110101010101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100111110101010101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100111110101010110) && ({row_reg, col_reg}<19'b0100111110111001011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100111110111001011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100111110111001100) && ({row_reg, col_reg}<19'b0100111110111001111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100111110111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100111110111010000) && ({row_reg, col_reg}<19'b0100111110111101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0100111110111101100) && ({row_reg, col_reg}<19'b0100111110111101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100111110111101110) && ({row_reg, col_reg}<19'b0100111111001110010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0100111111001110010) && ({row_reg, col_reg}<19'b0100111111001110100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0100111111001110100) && ({row_reg, col_reg}<19'b0100111111001110110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0100111111001110110) && ({row_reg, col_reg}<19'b0100111111001111000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0100111111001111000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100111111001111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0100111111001111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0100111111001111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0100111111001111100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0100111111001111101)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0100111111001111110) && ({row_reg, col_reg}<19'b0101000000010100011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101000000010100011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0101000000010100100)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=19'b0101000000010100101) && ({row_reg, col_reg}<19'b0101000001001111000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0101000001001111000) && ({row_reg, col_reg}<19'b0101000001001111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101000001001111010) && ({row_reg, col_reg}<19'b0101000001001111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101000001001111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101000001001111101)) color_data = 12'b101110111011;

		if(({row_reg, col_reg}>=19'b0101000001001111110) && ({row_reg, col_reg}<19'b0101000010010100010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101000010010100010)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0101000010010100011)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0101000010010100100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101000010010100101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101000010010100110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101000010010100111) && ({row_reg, col_reg}<19'b0101000011001111001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0101000011001111001) && ({row_reg, col_reg}<19'b0101000011001111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101000011001111011) && ({row_reg, col_reg}<19'b0101000011001111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101000011001111101)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0101000011001111110)) color_data = 12'b110111011101;

		if(({row_reg, col_reg}>=19'b0101000011001111111) && ({row_reg, col_reg}<19'b0101000100010100010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101000100010100010)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0101000100010100011)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=19'b0101000100010100100) && ({row_reg, col_reg}<19'b0101000100010100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101000100010100110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101000100010100111) && ({row_reg, col_reg}<19'b0101000101001111001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0101000101001111001) && ({row_reg, col_reg}<19'b0101000101001111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101000101001111011) && ({row_reg, col_reg}<19'b0101000101001111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101000101001111110)) color_data = 12'b101010101010;

		if(({row_reg, col_reg}==19'b0101000101001111111)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=19'b0101000110000000000) && ({row_reg, col_reg}<19'b0101000110010100001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101000110010100001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0101000110010100010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0101000110010100011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101000110010100100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101000110010100101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101000110010100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101000110010100111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101000110010101000) && ({row_reg, col_reg}<19'b0101000111001111000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101000111001111000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101000111001111001) && ({row_reg, col_reg}<19'b0101000111001111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101000111001111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101000111001111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101000111001111110)) color_data = 12'b100110011001;

		if(({row_reg, col_reg}==19'b0101000111001111111)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0101001000000000000) && ({row_reg, col_reg}<19'b0101001000010100001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101001000010100001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0101001000010100010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0101001000010100011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101001000010100100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101001000010100101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101001000010100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101001000010100111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101001000010101000) && ({row_reg, col_reg}<19'b0101001001001111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101001001001111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101001001001111011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101001001001111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101001001001111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101001001001111110)) color_data = 12'b100010001000;

		if(({row_reg, col_reg}==19'b0101001001001111111)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=19'b0101001010000000000) && ({row_reg, col_reg}<19'b0101001010010100001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101001010010100001)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0101001010010100010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=19'b0101001010010100011) && ({row_reg, col_reg}<19'b0101001010010100101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101001010010100101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101001010010100110) && ({row_reg, col_reg}<19'b0101001011001111000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101001011001111000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101001011001111001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101001011001111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101001011001111011) && ({row_reg, col_reg}<19'b0101001011001111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101001011001111110)) color_data = 12'b100010001000;

		if(({row_reg, col_reg}==19'b0101001011001111111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=19'b0101001100000000000) && ({row_reg, col_reg}<19'b0101001100010100001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101001100010100001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0101001100010100010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101001100010100011) && ({row_reg, col_reg}<19'b0101001100010100101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101001100010100101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101001100010100110) && ({row_reg, col_reg}<19'b0101001101001111000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101001101001111000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101001101001111001) && ({row_reg, col_reg}<19'b0101001101001111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0101001101001111101) && ({row_reg, col_reg}<19'b0101001101001111111)) color_data = 12'b100010001000;

		if(({row_reg, col_reg}==19'b0101001101001111111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=19'b0101001110000000000) && ({row_reg, col_reg}<19'b0101001110010100001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101001110010100001)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=19'b0101001110010100010) && ({row_reg, col_reg}<19'b0101001110010100100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101001110010100100) && ({row_reg, col_reg}<19'b0101001110010100111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101001110010100111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101001110010101000) && ({row_reg, col_reg}<19'b0101001111001111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0101001111001111010) && ({row_reg, col_reg}<19'b0101001111001111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101001111001111100) && ({row_reg, col_reg}<19'b0101001111001111111)) color_data = 12'b011101110111;

		if(({row_reg, col_reg}==19'b0101001111001111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101010000000000000) && ({row_reg, col_reg}<19'b0101010000010100001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101010000010100001)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0101010000010100010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101010000010100011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101010000010100100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101010000010100101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101010000010100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101010000010100111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101010000010101000) && ({row_reg, col_reg}<19'b0101010001001111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101010001001111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101010001001111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101010001001111110)) color_data = 12'b100010001000;

		if(({row_reg, col_reg}==19'b0101010001001111111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=19'b0101010010000000000) && ({row_reg, col_reg}<19'b0101010010010100001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101010010010100001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=19'b0101010010010100010) && ({row_reg, col_reg}<19'b0101010010010100100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101010010010100100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101010010010100101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101010010010100110) && ({row_reg, col_reg}<19'b0101010011001111000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0101010011001111000) && ({row_reg, col_reg}<19'b0101010011001111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101010011001111011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101010011001111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101010011001111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101010011001111110)) color_data = 12'b100010001000;

		if(({row_reg, col_reg}==19'b0101010011001111111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=19'b0101010100000000000) && ({row_reg, col_reg}<19'b0101010100010100001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101010100010100001)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0101010100010100010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0101010100010100011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0101010100010100100) && ({row_reg, col_reg}<19'b0101010100010100110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101010100010100110) && ({row_reg, col_reg}<19'b0101010101001111000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101010101001111000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101010101001111001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101010101001111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101010101001111011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101010101001111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101010101001111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101010101001111110)) color_data = 12'b100010001000;

		if(({row_reg, col_reg}==19'b0101010101001111111)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=19'b0101010110000000000) && ({row_reg, col_reg}<19'b0101010110010100001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101010110010100001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0101010110010100010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0101010110010100011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0101010110010100100) && ({row_reg, col_reg}<19'b0101010110010100110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101010110010100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101010110010100111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101010110010101000) && ({row_reg, col_reg}<19'b0101010111001111000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101010111001111000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101010111001111001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101010111001111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101010111001111011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101010111001111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101010111001111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101010111001111110)) color_data = 12'b100010001000;

		if(({row_reg, col_reg}==19'b0101010111001111111)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=19'b0101011000000000000) && ({row_reg, col_reg}<19'b0101011000010100010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101011000010100010)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0101011000010100011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101011000010100100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101011000010100101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101011000010100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101011000010100111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101011000010101000) && ({row_reg, col_reg}<19'b0101011001001111000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101011001001111000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101011001001111001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0101011001001111010) && ({row_reg, col_reg}<19'b0101011001001111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101011001001111100) && ({row_reg, col_reg}<19'b0101011001001111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101011001001111110)) color_data = 12'b100110011001;

		if(({row_reg, col_reg}==19'b0101011001001111111)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0101011010000000000) && ({row_reg, col_reg}<19'b0101011010010100010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101011010010100010)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0101011010010100011)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=19'b0101011010010100100) && ({row_reg, col_reg}<19'b0101011011001111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0101011011001111010) && ({row_reg, col_reg}<19'b0101011011001111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101011011001111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101011011001111101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101011011001111110)) color_data = 12'b101110111011;

		if(({row_reg, col_reg}==19'b0101011011001111111)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=19'b0101011100000000000) && ({row_reg, col_reg}<19'b0101011100010100010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101011100010100010)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0101011100010100011)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0101011100010100100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101011100010100101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101011100010100110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101011100010100111) && ({row_reg, col_reg}<19'b0101011101001111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101011101001111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101011101001111101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0101011101001111110)) color_data = 12'b110111011101;

		if(({row_reg, col_reg}>=19'b0101011101001111111) && ({row_reg, col_reg}<19'b0101011110010100011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101011110010100011)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0101011110010100100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=19'b0101011110010100101) && ({row_reg, col_reg}<19'b0101011110010100111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101011110010100111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101011110010101000) && ({row_reg, col_reg}<19'b0101011111001111000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0101011111001111000) && ({row_reg, col_reg}<19'b0101011111001111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101011111001111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0101011111001111011) && ({row_reg, col_reg}<19'b0101011111001111101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101011111001111101)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=19'b0101011111001111110) && ({row_reg, col_reg}<19'b0101100000010100100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101100000010100100)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0101100000010100101)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=19'b0101100000010100110) && ({row_reg, col_reg}<19'b0101100000010101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0101100000010101101) && ({row_reg, col_reg}<19'b0101100000010101111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101100000010101111) && ({row_reg, col_reg}<19'b0101100000100111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101100000100111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101100000100111011) && ({row_reg, col_reg}<19'b0101100000100111111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101100000100111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101100000101000000) && ({row_reg, col_reg}<19'b0101100000101010000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101100000101010000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101100000101010001) && ({row_reg, col_reg}<19'b0101100000101010100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101100000101010100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101100000101010101) && ({row_reg, col_reg}<19'b0101100000101010111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101100000101010111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101100000101011000) && ({row_reg, col_reg}<19'b0101100000111001000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101100000111001000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101100000111001001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101100000111001010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101100000111001011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101100000111001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101100000111001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101100000111001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101100000111001111) && ({row_reg, col_reg}<19'b0101100000111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0101100000111101000) && ({row_reg, col_reg}<19'b0101100000111101010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101100000111101010) && ({row_reg, col_reg}<19'b0101100000111101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101100000111101101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101100000111101110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101100000111101111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101100000111110000) && ({row_reg, col_reg}<19'b0101100001001110000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0101100001001110000) && ({row_reg, col_reg}<19'b0101100001001110010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101100001001110010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0101100001001110011) && ({row_reg, col_reg}<19'b0101100001001110110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101100001001110110) && ({row_reg, col_reg}<19'b0101100001001111000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101100001001111000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101100001001111001) && ({row_reg, col_reg}<19'b0101100001001111011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101100001001111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101100001001111100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0101100001001111101)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0101100001001111110) && ({row_reg, col_reg}<19'b0101100010010100100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101100010010100100)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0101100010010100101)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0101100010010100110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0101100010010100111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101100010010101000) && ({row_reg, col_reg}<19'b0101100010010101010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0101100010010101010) && ({row_reg, col_reg}<19'b0101100010010101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101100010010101100) && ({row_reg, col_reg}<19'b0101100010100111000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101100010100111000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101100010100111001) && ({row_reg, col_reg}<19'b0101100010101010010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101100010101010010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101100010101010011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0101100010101010100) && ({row_reg, col_reg}<19'b0101100010101010110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101100010101010110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101100010101010111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101100010101011000) && ({row_reg, col_reg}<19'b0101100010111001010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101100010111001010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101100010111001011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0101100010111001100) && ({row_reg, col_reg}<19'b0101100010111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101100010111001111) && ({row_reg, col_reg}<19'b0101100010111101001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0101100010111101001) && ({row_reg, col_reg}<19'b0101100010111101011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101100010111101011) && ({row_reg, col_reg}<19'b0101100010111101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101100010111101101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101100010111101110) && ({row_reg, col_reg}<19'b0101100011001110000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101100011001110000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101100011001110001) && ({row_reg, col_reg}<19'b0101100011001110101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0101100011001110101) && ({row_reg, col_reg}<19'b0101100011001111000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101100011001111000) && ({row_reg, col_reg}<19'b0101100011001111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101100011001111010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0101100011001111011)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0101100011001111100)) color_data = 12'b110111011101;

		if(({row_reg, col_reg}>=19'b0101100011001111101) && ({row_reg, col_reg}<19'b0101100100010100110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101100100010100110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0101100100010100111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=19'b0101100100010101000) && ({row_reg, col_reg}<19'b0101100100010101010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101100100010101010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0101100100010101011) && ({row_reg, col_reg}<19'b0101100100100111000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101100100100111000) && ({row_reg, col_reg}<19'b0101100100100111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101100100100111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101100100100111011) && ({row_reg, col_reg}<19'b0101100100100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101100100100111101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101100100100111110) && ({row_reg, col_reg}<19'b0101100100101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0101100100101010001) && ({row_reg, col_reg}<19'b0101100100101010011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101100100101010011) && ({row_reg, col_reg}<19'b0101100100101011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0101100100101011000) && ({row_reg, col_reg}<19'b0101100100111001001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101100100111001001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101100100111001010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101100100111001011) && ({row_reg, col_reg}<19'b0101100100111101001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0101100100111101001) && ({row_reg, col_reg}<19'b0101100100111101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101100100111101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0101100100111101101) && ({row_reg, col_reg}<19'b0101100100111101111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101100100111101111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0101100100111110000) && ({row_reg, col_reg}<19'b0101100101001110000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101100101001110000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0101100101001110001) && ({row_reg, col_reg}<19'b0101100101001110101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101100101001110101) && ({row_reg, col_reg}<19'b0101100101001111000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101100101001111000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101100101001111001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0101100101001111010)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0101100101001111011)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0101100101001111100) && ({row_reg, col_reg}<19'b0101100110010100111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101100110010100111)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0101100110010101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0101100110010101001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=19'b0101100110010101010) && ({row_reg, col_reg}<19'b0101100110010101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101100110010101100) && ({row_reg, col_reg}<19'b0101100110100111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101100110100111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101100110100111011) && ({row_reg, col_reg}<19'b0101100110100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101100110100111101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101100110100111110) && ({row_reg, col_reg}<19'b0101100110101010101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0101100110101010101) && ({row_reg, col_reg}<19'b0101100110101011000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101100110101011000) && ({row_reg, col_reg}<19'b0101100110111001010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101100110111001010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101100110111001011) && ({row_reg, col_reg}<19'b0101100110111001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0101100110111001101) && ({row_reg, col_reg}<19'b0101100110111010000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101100110111010000) && ({row_reg, col_reg}<19'b0101100110111101001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101100110111101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101100110111101010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101100110111101011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101100110111101100) && ({row_reg, col_reg}<19'b0101100111001110101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0101100111001110101) && ({row_reg, col_reg}<19'b0101100111001110111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101100111001110111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0101100111001111000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0101100111001111001)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0101100111001111010)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0101100111001111011) && ({row_reg, col_reg}<19'b0101101000010101001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101101000010101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b0101101000010101010)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=19'b0101101000010101011) && ({row_reg, col_reg}<19'b0101101000010101101)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0101101000010101101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=19'b0101101000010101110) && ({row_reg, col_reg}<19'b0101101000100111001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=19'b0101101000100111001) && ({row_reg, col_reg}<19'b0101101000100111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101101000100111011) && ({row_reg, col_reg}<19'b0101101000100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101101000100111101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101101000100111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101101000100111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101101000101000000) && ({row_reg, col_reg}<19'b0101101000101010000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b0101101000101010000) && ({row_reg, col_reg}<19'b0101101000101010011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101101000101010011) && ({row_reg, col_reg}<19'b0101101000111001110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0101101000111001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101101000111001111) && ({row_reg, col_reg}<19'b0101101000111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101101000111101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101101000111101001) && ({row_reg, col_reg}<19'b0101101001001110100)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0101101001001110100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0101101001001110101)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0101101001001110110)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0101101001001110111)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0101101001001111000)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0101101001001111001) && ({row_reg, col_reg}<19'b0101101010010101101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101101010010101101)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=19'b0101101010010101110) && ({row_reg, col_reg}<19'b0101101010100111000)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0101101010100111000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0101101010100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101101010100111010) && ({row_reg, col_reg}<19'b0101101010100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101101010100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101101010100111101) && ({row_reg, col_reg}<19'b0101101010100111111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101101010100111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101101010101000000) && ({row_reg, col_reg}<19'b0101101010101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101101010101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101101010101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0101101010101010011)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=19'b0101101010101010100) && ({row_reg, col_reg}<19'b0101101010101010111)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0101101010101010111)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=19'b0101101010101011000) && ({row_reg, col_reg}<19'b0101101010111001000)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0101101010111001000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=19'b0101101010111001001) && ({row_reg, col_reg}<19'b0101101010111001110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0101101010111001110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0101101010111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101101010111010000) && ({row_reg, col_reg}<19'b0101101010111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101101010111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=19'b0101101010111101001) && ({row_reg, col_reg}<19'b0101101011001110011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0101101011001110011) && ({row_reg, col_reg}<19'b0101101011001110101)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0101101011001110101) && ({row_reg, col_reg}<19'b0101101100100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101101100100111000)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b0101101100100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101101100100111010) && ({row_reg, col_reg}<19'b0101101100100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101101100100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101101100100111101) && ({row_reg, col_reg}<19'b0101101100100111111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101101100100111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101101100101000000) && ({row_reg, col_reg}<19'b0101101100101010010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101101100101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0101101100101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0101101100101010100) && ({row_reg, col_reg}<19'b0101101100111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101101100111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0101101100111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101101100111010000) && ({row_reg, col_reg}<19'b0101101100111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101101100111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0101101100111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0101101100111101010) && ({row_reg, col_reg}<19'b0101101110100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101101110100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=19'b0101101110100111001) && ({row_reg, col_reg}<19'b0101101110100111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101101110100111011) && ({row_reg, col_reg}<19'b0101101110100111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101101110100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101101110100111111) && ({row_reg, col_reg}<19'b0101101110101010000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101101110101010000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101101110101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101101110101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0101101110101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0101101110101010100) && ({row_reg, col_reg}<19'b0101101110111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101101110111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0101101110111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101101110111010000) && ({row_reg, col_reg}<19'b0101101110111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101101110111101000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0101101110111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0101101110111101010) && ({row_reg, col_reg}<19'b0101110000100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101110000100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0101110000100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101110000100111010) && ({row_reg, col_reg}<19'b0101110000100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101110000100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101110000100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101110000100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101110000100111111) && ({row_reg, col_reg}<19'b0101110000101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101110000101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101110000101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0101110000101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0101110000101010100) && ({row_reg, col_reg}<19'b0101110000111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101110000111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0101110000111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101110000111010000) && ({row_reg, col_reg}<19'b0101110000111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101110000111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0101110000111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0101110000111101010) && ({row_reg, col_reg}<19'b0101110010100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101110010100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0101110010100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101110010100111010) && ({row_reg, col_reg}<19'b0101110010100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101110010100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101110010100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101110010100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101110010100111111) && ({row_reg, col_reg}<19'b0101110010101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101110010101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101110010101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0101110010101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0101110010101010100) && ({row_reg, col_reg}<19'b0101110010111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101110010111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0101110010111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101110010111010000) && ({row_reg, col_reg}<19'b0101110010111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101110010111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0101110010111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0101110010111101010) && ({row_reg, col_reg}<19'b0101110100100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101110100100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0101110100100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101110100100111010) && ({row_reg, col_reg}<19'b0101110100100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101110100100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101110100100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101110100100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101110100100111111) && ({row_reg, col_reg}<19'b0101110100101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101110100101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101110100101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0101110100101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0101110100101010100) && ({row_reg, col_reg}<19'b0101110100111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101110100111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0101110100111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101110100111010000) && ({row_reg, col_reg}<19'b0101110100111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101110100111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0101110100111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0101110100111101010) && ({row_reg, col_reg}<19'b0101110110100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101110110100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0101110110100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101110110100111010) && ({row_reg, col_reg}<19'b0101110110100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101110110100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101110110100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101110110100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101110110100111111) && ({row_reg, col_reg}<19'b0101110110101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101110110101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101110110101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0101110110101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0101110110101010100) && ({row_reg, col_reg}<19'b0101110110111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101110110111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0101110110111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101110110111010000) && ({row_reg, col_reg}<19'b0101110110111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101110110111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0101110110111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0101110110111101010) && ({row_reg, col_reg}<19'b0101111000100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101111000100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0101111000100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101111000100111010) && ({row_reg, col_reg}<19'b0101111000100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101111000100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101111000100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101111000100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101111000100111111) && ({row_reg, col_reg}<19'b0101111000101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101111000101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101111000101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0101111000101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0101111000101010100) && ({row_reg, col_reg}<19'b0101111000111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101111000111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0101111000111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101111000111010000) && ({row_reg, col_reg}<19'b0101111000111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101111000111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0101111000111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0101111000111101010) && ({row_reg, col_reg}<19'b0101111010100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101111010100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0101111010100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101111010100111010) && ({row_reg, col_reg}<19'b0101111010100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101111010100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101111010100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101111010100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101111010100111111) && ({row_reg, col_reg}<19'b0101111010101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101111010101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101111010101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0101111010101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0101111010101010100) && ({row_reg, col_reg}<19'b0101111010111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101111010111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0101111010111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101111010111010000) && ({row_reg, col_reg}<19'b0101111010111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101111010111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0101111010111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0101111010111101010) && ({row_reg, col_reg}<19'b0101111100100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101111100100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0101111100100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101111100100111010) && ({row_reg, col_reg}<19'b0101111100100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101111100100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101111100100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101111100100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101111100100111111) && ({row_reg, col_reg}<19'b0101111100101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101111100101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101111100101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0101111100101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0101111100101010100) && ({row_reg, col_reg}<19'b0101111100111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101111100111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0101111100111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101111100111010000) && ({row_reg, col_reg}<19'b0101111100111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101111100111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0101111100111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0101111100111101010) && ({row_reg, col_reg}<19'b0101111110100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101111110100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0101111110100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101111110100111010) && ({row_reg, col_reg}<19'b0101111110100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101111110100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101111110100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101111110100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101111110100111111) && ({row_reg, col_reg}<19'b0101111110101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101111110101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0101111110101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0101111110101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0101111110101010100) && ({row_reg, col_reg}<19'b0101111110111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0101111110111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0101111110111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0101111110111010000) && ({row_reg, col_reg}<19'b0101111110111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0101111110111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0101111110111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0101111110111101010) && ({row_reg, col_reg}<19'b0110000000100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0110000000100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0110000000100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0110000000100111010) && ({row_reg, col_reg}<19'b0110000000100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110000000100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0110000000100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110000000100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0110000000100111111) && ({row_reg, col_reg}<19'b0110000000101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110000000101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0110000000101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0110000000101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0110000000101010100) && ({row_reg, col_reg}<19'b0110000000111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0110000000111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0110000000111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0110000000111010000) && ({row_reg, col_reg}<19'b0110000000111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110000000111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0110000000111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0110000000111101010) && ({row_reg, col_reg}<19'b0110000010100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0110000010100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0110000010100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0110000010100111010) && ({row_reg, col_reg}<19'b0110000010100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110000010100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0110000010100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110000010100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0110000010100111111) && ({row_reg, col_reg}<19'b0110000010101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110000010101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0110000010101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0110000010101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0110000010101010100) && ({row_reg, col_reg}<19'b0110000010111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0110000010111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0110000010111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0110000010111010000) && ({row_reg, col_reg}<19'b0110000010111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110000010111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0110000010111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0110000010111101010) && ({row_reg, col_reg}<19'b0110000100100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0110000100100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0110000100100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0110000100100111010) && ({row_reg, col_reg}<19'b0110000100100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110000100100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0110000100100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110000100100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0110000100100111111) && ({row_reg, col_reg}<19'b0110000100101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110000100101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0110000100101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0110000100101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0110000100101010100) && ({row_reg, col_reg}<19'b0110000100111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0110000100111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0110000100111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0110000100111010000) && ({row_reg, col_reg}<19'b0110000100111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110000100111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0110000100111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0110000100111101010) && ({row_reg, col_reg}<19'b0110000110100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0110000110100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0110000110100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0110000110100111010) && ({row_reg, col_reg}<19'b0110000110100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110000110100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0110000110100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110000110100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0110000110100111111) && ({row_reg, col_reg}<19'b0110000110101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110000110101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0110000110101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0110000110101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0110000110101010100) && ({row_reg, col_reg}<19'b0110000110111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0110000110111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0110000110111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0110000110111010000) && ({row_reg, col_reg}<19'b0110000110111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110000110111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0110000110111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0110000110111101010) && ({row_reg, col_reg}<19'b0110001000100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0110001000100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0110001000100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0110001000100111010) && ({row_reg, col_reg}<19'b0110001000100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110001000100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0110001000100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110001000100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0110001000100111111) && ({row_reg, col_reg}<19'b0110001000101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110001000101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0110001000101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0110001000101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0110001000101010100) && ({row_reg, col_reg}<19'b0110001000111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0110001000111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0110001000111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0110001000111010000) && ({row_reg, col_reg}<19'b0110001000111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110001000111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0110001000111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0110001000111101010) && ({row_reg, col_reg}<19'b0110001010100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0110001010100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0110001010100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0110001010100111010) && ({row_reg, col_reg}<19'b0110001010100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110001010100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0110001010100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110001010100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0110001010100111111) && ({row_reg, col_reg}<19'b0110001010101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110001010101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0110001010101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0110001010101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0110001010101010100) && ({row_reg, col_reg}<19'b0110001010111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0110001010111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0110001010111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0110001010111010000) && ({row_reg, col_reg}<19'b0110001010111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110001010111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0110001010111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0110001010111101010) && ({row_reg, col_reg}<19'b0110001100100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0110001100100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0110001100100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0110001100100111010) && ({row_reg, col_reg}<19'b0110001100100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110001100100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0110001100100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110001100100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0110001100100111111) && ({row_reg, col_reg}<19'b0110001100101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110001100101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0110001100101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0110001100101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0110001100101010100) && ({row_reg, col_reg}<19'b0110001100111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0110001100111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0110001100111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0110001100111010000) && ({row_reg, col_reg}<19'b0110001100111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110001100111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0110001100111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0110001100111101010) && ({row_reg, col_reg}<19'b0110001110100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0110001110100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0110001110100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0110001110100111010) && ({row_reg, col_reg}<19'b0110001110100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110001110100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0110001110100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110001110100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0110001110100111111) && ({row_reg, col_reg}<19'b0110001110101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110001110101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0110001110101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0110001110101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0110001110101010100) && ({row_reg, col_reg}<19'b0110001110111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0110001110111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0110001110111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0110001110111010000) && ({row_reg, col_reg}<19'b0110001110111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110001110111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0110001110111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0110001110111101010) && ({row_reg, col_reg}<19'b0110010000100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0110010000100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0110010000100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0110010000100111010) && ({row_reg, col_reg}<19'b0110010000100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110010000100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0110010000100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110010000100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0110010000100111111) && ({row_reg, col_reg}<19'b0110010000101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110010000101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0110010000101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0110010000101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0110010000101010100) && ({row_reg, col_reg}<19'b0110010000111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0110010000111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0110010000111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0110010000111010000) && ({row_reg, col_reg}<19'b0110010000111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110010000111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0110010000111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0110010000111101010) && ({row_reg, col_reg}<19'b0110010010100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0110010010100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0110010010100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0110010010100111010) && ({row_reg, col_reg}<19'b0110010010100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110010010100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0110010010100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110010010100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0110010010100111111) && ({row_reg, col_reg}<19'b0110010010101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110010010101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0110010010101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0110010010101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0110010010101010100) && ({row_reg, col_reg}<19'b0110010010111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0110010010111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0110010010111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0110010010111010000) && ({row_reg, col_reg}<19'b0110010010111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110010010111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0110010010111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0110010010111101010) && ({row_reg, col_reg}<19'b0110010100100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0110010100100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0110010100100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0110010100100111010) && ({row_reg, col_reg}<19'b0110010100100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110010100100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0110010100100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110010100100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0110010100100111111) && ({row_reg, col_reg}<19'b0110010100101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110010100101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0110010100101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0110010100101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0110010100101010100) && ({row_reg, col_reg}<19'b0110010100111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0110010100111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0110010100111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0110010100111010000) && ({row_reg, col_reg}<19'b0110010100111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110010100111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0110010100111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0110010100111101010) && ({row_reg, col_reg}<19'b0110010110100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0110010110100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0110010110100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0110010110100111010) && ({row_reg, col_reg}<19'b0110010110100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110010110100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0110010110100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110010110100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0110010110100111111) && ({row_reg, col_reg}<19'b0110010110101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110010110101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0110010110101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0110010110101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0110010110101010100) && ({row_reg, col_reg}<19'b0110010110111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0110010110111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0110010110111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0110010110111010000) && ({row_reg, col_reg}<19'b0110010110111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110010110111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0110010110111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0110010110111101010) && ({row_reg, col_reg}<19'b0110011000100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0110011000100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0110011000100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0110011000100111010) && ({row_reg, col_reg}<19'b0110011000100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110011000100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0110011000100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110011000100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0110011000100111111) && ({row_reg, col_reg}<19'b0110011000101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110011000101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0110011000101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0110011000101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0110011000101010100) && ({row_reg, col_reg}<19'b0110011000111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0110011000111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0110011000111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0110011000111010000) && ({row_reg, col_reg}<19'b0110011000111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110011000111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0110011000111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0110011000111101010) && ({row_reg, col_reg}<19'b0110011010100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0110011010100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0110011010100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0110011010100111010) && ({row_reg, col_reg}<19'b0110011010100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110011010100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0110011010100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110011010100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0110011010100111111) && ({row_reg, col_reg}<19'b0110011010101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110011010101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0110011010101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0110011010101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0110011010101010100) && ({row_reg, col_reg}<19'b0110011010111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0110011010111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0110011010111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0110011010111010000) && ({row_reg, col_reg}<19'b0110011010111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110011010111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0110011010111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0110011010111101010) && ({row_reg, col_reg}<19'b0110011100100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0110011100100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0110011100100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0110011100100111010) && ({row_reg, col_reg}<19'b0110011100100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110011100100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0110011100100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110011100100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0110011100100111111) && ({row_reg, col_reg}<19'b0110011100101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110011100101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0110011100101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0110011100101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0110011100101010100) && ({row_reg, col_reg}<19'b0110011100111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0110011100111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0110011100111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0110011100111010000) && ({row_reg, col_reg}<19'b0110011100111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110011100111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0110011100111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0110011100111101010) && ({row_reg, col_reg}<19'b0110011110100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0110011110100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0110011110100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0110011110100111010) && ({row_reg, col_reg}<19'b0110011110100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110011110100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0110011110100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110011110100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0110011110100111111) && ({row_reg, col_reg}<19'b0110011110101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110011110101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0110011110101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0110011110101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0110011110101010100) && ({row_reg, col_reg}<19'b0110011110111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0110011110111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0110011110111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0110011110111010000) && ({row_reg, col_reg}<19'b0110011110111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110011110111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0110011110111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0110011110111101010) && ({row_reg, col_reg}<19'b0110100000100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0110100000100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0110100000100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0110100000100111010) && ({row_reg, col_reg}<19'b0110100000100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110100000100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0110100000100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110100000100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0110100000100111111) && ({row_reg, col_reg}<19'b0110100000101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110100000101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0110100000101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0110100000101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0110100000101010100) && ({row_reg, col_reg}<19'b0110100000111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0110100000111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0110100000111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0110100000111010000) && ({row_reg, col_reg}<19'b0110100000111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110100000111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0110100000111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0110100000111101010) && ({row_reg, col_reg}<19'b0110100010100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0110100010100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0110100010100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0110100010100111010) && ({row_reg, col_reg}<19'b0110100010100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110100010100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0110100010100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110100010100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0110100010100111111) && ({row_reg, col_reg}<19'b0110100010101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110100010101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0110100010101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0110100010101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0110100010101010100) && ({row_reg, col_reg}<19'b0110100010111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0110100010111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0110100010111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0110100010111010000) && ({row_reg, col_reg}<19'b0110100010111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110100010111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0110100010111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0110100010111101010) && ({row_reg, col_reg}<19'b0110100100100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0110100100100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0110100100100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0110100100100111010) && ({row_reg, col_reg}<19'b0110100100100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110100100100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0110100100100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110100100100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0110100100100111111) && ({row_reg, col_reg}<19'b0110100100101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110100100101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0110100100101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0110100100101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0110100100101010100) && ({row_reg, col_reg}<19'b0110100100111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0110100100111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0110100100111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0110100100111010000) && ({row_reg, col_reg}<19'b0110100100111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110100100111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0110100100111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0110100100111101010) && ({row_reg, col_reg}<19'b0110100110100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0110100110100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0110100110100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0110100110100111010) && ({row_reg, col_reg}<19'b0110100110100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110100110100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0110100110100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110100110100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0110100110100111111) && ({row_reg, col_reg}<19'b0110100110101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110100110101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0110100110101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0110100110101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0110100110101010100) && ({row_reg, col_reg}<19'b0110100110111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0110100110111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0110100110111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0110100110111010000) && ({row_reg, col_reg}<19'b0110100110111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110100110111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0110100110111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0110100110111101010) && ({row_reg, col_reg}<19'b0110101000100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0110101000100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0110101000100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0110101000100111010) && ({row_reg, col_reg}<19'b0110101000100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110101000100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0110101000100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110101000100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0110101000100111111) && ({row_reg, col_reg}<19'b0110101000101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110101000101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0110101000101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0110101000101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0110101000101010100) && ({row_reg, col_reg}<19'b0110101000111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0110101000111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0110101000111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0110101000111010000) && ({row_reg, col_reg}<19'b0110101000111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110101000111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0110101000111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0110101000111101010) && ({row_reg, col_reg}<19'b0110101010100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0110101010100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0110101010100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0110101010100111010) && ({row_reg, col_reg}<19'b0110101010100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110101010100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0110101010100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110101010100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0110101010100111111) && ({row_reg, col_reg}<19'b0110101010101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110101010101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0110101010101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0110101010101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0110101010101010100) && ({row_reg, col_reg}<19'b0110101010111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0110101010111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0110101010111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0110101010111010000) && ({row_reg, col_reg}<19'b0110101010111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110101010111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0110101010111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0110101010111101010) && ({row_reg, col_reg}<19'b0110101100100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0110101100100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0110101100100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0110101100100111010) && ({row_reg, col_reg}<19'b0110101100100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110101100100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0110101100100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110101100100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0110101100100111111) && ({row_reg, col_reg}<19'b0110101100101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110101100101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0110101100101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0110101100101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0110101100101010100) && ({row_reg, col_reg}<19'b0110101100111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0110101100111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0110101100111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0110101100111010000) && ({row_reg, col_reg}<19'b0110101100111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110101100111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0110101100111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0110101100111101010) && ({row_reg, col_reg}<19'b0110101110100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0110101110100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0110101110100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0110101110100111010) && ({row_reg, col_reg}<19'b0110101110100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110101110100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0110101110100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110101110100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0110101110100111111) && ({row_reg, col_reg}<19'b0110101110101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110101110101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0110101110101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0110101110101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0110101110101010100) && ({row_reg, col_reg}<19'b0110101110111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0110101110111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0110101110111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0110101110111010000) && ({row_reg, col_reg}<19'b0110101110111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110101110111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0110101110111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0110101110111101010) && ({row_reg, col_reg}<19'b0110110000100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0110110000100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0110110000100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0110110000100111010) && ({row_reg, col_reg}<19'b0110110000100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110110000100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0110110000100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110110000100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0110110000100111111) && ({row_reg, col_reg}<19'b0110110000101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110110000101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0110110000101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0110110000101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0110110000101010100) && ({row_reg, col_reg}<19'b0110110000111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0110110000111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0110110000111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0110110000111010000) && ({row_reg, col_reg}<19'b0110110000111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110110000111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0110110000111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0110110000111101010) && ({row_reg, col_reg}<19'b0110110010100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0110110010100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0110110010100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0110110010100111010) && ({row_reg, col_reg}<19'b0110110010100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110110010100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0110110010100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110110010100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0110110010100111111) && ({row_reg, col_reg}<19'b0110110010101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110110010101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0110110010101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0110110010101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0110110010101010100) && ({row_reg, col_reg}<19'b0110110010111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0110110010111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0110110010111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0110110010111010000) && ({row_reg, col_reg}<19'b0110110010111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110110010111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0110110010111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0110110010111101010) && ({row_reg, col_reg}<19'b0110110100100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0110110100100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0110110100100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0110110100100111010) && ({row_reg, col_reg}<19'b0110110100100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110110100100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0110110100100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110110100100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0110110100100111111) && ({row_reg, col_reg}<19'b0110110100101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110110100101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0110110100101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0110110100101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0110110100101010100) && ({row_reg, col_reg}<19'b0110110100111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0110110100111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0110110100111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0110110100111010000) && ({row_reg, col_reg}<19'b0110110100111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110110100111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0110110100111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0110110100111101010) && ({row_reg, col_reg}<19'b0110110110100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0110110110100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0110110110100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0110110110100111010) && ({row_reg, col_reg}<19'b0110110110100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110110110100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0110110110100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110110110100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0110110110100111111) && ({row_reg, col_reg}<19'b0110110110101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110110110101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0110110110101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0110110110101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0110110110101010100) && ({row_reg, col_reg}<19'b0110110110111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0110110110111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0110110110111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0110110110111010000) && ({row_reg, col_reg}<19'b0110110110111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110110110111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0110110110111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0110110110111101010) && ({row_reg, col_reg}<19'b0110111000100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0110111000100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0110111000100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0110111000100111010) && ({row_reg, col_reg}<19'b0110111000100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110111000100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0110111000100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110111000100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0110111000100111111) && ({row_reg, col_reg}<19'b0110111000101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110111000101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0110111000101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0110111000101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0110111000101010100) && ({row_reg, col_reg}<19'b0110111000111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0110111000111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0110111000111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0110111000111010000) && ({row_reg, col_reg}<19'b0110111000111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110111000111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0110111000111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0110111000111101010) && ({row_reg, col_reg}<19'b0110111010100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0110111010100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0110111010100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0110111010100111010) && ({row_reg, col_reg}<19'b0110111010100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110111010100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0110111010100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110111010100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0110111010100111111) && ({row_reg, col_reg}<19'b0110111010101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110111010101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0110111010101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0110111010101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0110111010101010100) && ({row_reg, col_reg}<19'b0110111010111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0110111010111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0110111010111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0110111010111010000) && ({row_reg, col_reg}<19'b0110111010111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110111010111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0110111010111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0110111010111101010) && ({row_reg, col_reg}<19'b0110111100100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0110111100100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0110111100100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0110111100100111010) && ({row_reg, col_reg}<19'b0110111100100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110111100100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0110111100100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110111100100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0110111100100111111) && ({row_reg, col_reg}<19'b0110111100101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110111100101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0110111100101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0110111100101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0110111100101010100) && ({row_reg, col_reg}<19'b0110111100111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0110111100111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0110111100111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0110111100111010000) && ({row_reg, col_reg}<19'b0110111100111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110111100111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0110111100111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0110111100111101010) && ({row_reg, col_reg}<19'b0110111110100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0110111110100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0110111110100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0110111110100111010) && ({row_reg, col_reg}<19'b0110111110100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110111110100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0110111110100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110111110100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0110111110100111111) && ({row_reg, col_reg}<19'b0110111110101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110111110101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0110111110101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0110111110101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0110111110101010100) && ({row_reg, col_reg}<19'b0110111110111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0110111110111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0110111110111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0110111110111010000) && ({row_reg, col_reg}<19'b0110111110111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0110111110111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0110111110111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0110111110111101010) && ({row_reg, col_reg}<19'b0111000000100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111000000100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0111000000100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111000000100111010) && ({row_reg, col_reg}<19'b0111000000100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111000000100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0111000000100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111000000100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111000000100111111) && ({row_reg, col_reg}<19'b0111000000101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111000000101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0111000000101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0111000000101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0111000000101010100) && ({row_reg, col_reg}<19'b0111000000111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111000000111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0111000000111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111000000111010000) && ({row_reg, col_reg}<19'b0111000000111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111000000111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0111000000111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0111000000111101010) && ({row_reg, col_reg}<19'b0111000010100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111000010100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0111000010100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111000010100111010) && ({row_reg, col_reg}<19'b0111000010100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111000010100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0111000010100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111000010100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111000010100111111) && ({row_reg, col_reg}<19'b0111000010101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111000010101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0111000010101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0111000010101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0111000010101010100) && ({row_reg, col_reg}<19'b0111000010111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111000010111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0111000010111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111000010111010000) && ({row_reg, col_reg}<19'b0111000010111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111000010111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0111000010111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0111000010111101010) && ({row_reg, col_reg}<19'b0111000100100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111000100100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0111000100100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111000100100111010) && ({row_reg, col_reg}<19'b0111000100100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111000100100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0111000100100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111000100100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111000100100111111) && ({row_reg, col_reg}<19'b0111000100101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111000100101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0111000100101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0111000100101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0111000100101010100) && ({row_reg, col_reg}<19'b0111000100111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111000100111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0111000100111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111000100111010000) && ({row_reg, col_reg}<19'b0111000100111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111000100111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0111000100111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0111000100111101010) && ({row_reg, col_reg}<19'b0111000110100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111000110100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0111000110100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111000110100111010) && ({row_reg, col_reg}<19'b0111000110100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111000110100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0111000110100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111000110100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111000110100111111) && ({row_reg, col_reg}<19'b0111000110101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111000110101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0111000110101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0111000110101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0111000110101010100) && ({row_reg, col_reg}<19'b0111000110111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111000110111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0111000110111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111000110111010000) && ({row_reg, col_reg}<19'b0111000110111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111000110111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0111000110111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0111000110111101010) && ({row_reg, col_reg}<19'b0111001000100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111001000100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0111001000100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111001000100111010) && ({row_reg, col_reg}<19'b0111001000100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111001000100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0111001000100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111001000100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111001000100111111) && ({row_reg, col_reg}<19'b0111001000101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111001000101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0111001000101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0111001000101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0111001000101010100) && ({row_reg, col_reg}<19'b0111001000111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111001000111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0111001000111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111001000111010000) && ({row_reg, col_reg}<19'b0111001000111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111001000111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0111001000111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0111001000111101010) && ({row_reg, col_reg}<19'b0111001010100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111001010100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0111001010100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111001010100111010) && ({row_reg, col_reg}<19'b0111001010100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111001010100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0111001010100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111001010100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111001010100111111) && ({row_reg, col_reg}<19'b0111001010101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111001010101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0111001010101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0111001010101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0111001010101010100) && ({row_reg, col_reg}<19'b0111001010111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111001010111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0111001010111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111001010111010000) && ({row_reg, col_reg}<19'b0111001010111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111001010111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0111001010111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0111001010111101010) && ({row_reg, col_reg}<19'b0111001100100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111001100100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0111001100100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111001100100111010) && ({row_reg, col_reg}<19'b0111001100100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111001100100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0111001100100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111001100100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111001100100111111) && ({row_reg, col_reg}<19'b0111001100101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111001100101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0111001100101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0111001100101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0111001100101010100) && ({row_reg, col_reg}<19'b0111001100111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111001100111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0111001100111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111001100111010000) && ({row_reg, col_reg}<19'b0111001100111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111001100111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0111001100111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0111001100111101010) && ({row_reg, col_reg}<19'b0111001110100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111001110100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0111001110100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111001110100111010) && ({row_reg, col_reg}<19'b0111001110100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111001110100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0111001110100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111001110100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111001110100111111) && ({row_reg, col_reg}<19'b0111001110101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111001110101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0111001110101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0111001110101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0111001110101010100) && ({row_reg, col_reg}<19'b0111001110111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111001110111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0111001110111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111001110111010000) && ({row_reg, col_reg}<19'b0111001110111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111001110111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0111001110111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0111001110111101010) && ({row_reg, col_reg}<19'b0111010000100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111010000100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0111010000100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111010000100111010) && ({row_reg, col_reg}<19'b0111010000100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111010000100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0111010000100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111010000100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111010000100111111) && ({row_reg, col_reg}<19'b0111010000101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111010000101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0111010000101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0111010000101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0111010000101010100) && ({row_reg, col_reg}<19'b0111010000111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111010000111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0111010000111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111010000111010000) && ({row_reg, col_reg}<19'b0111010000111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111010000111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0111010000111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0111010000111101010) && ({row_reg, col_reg}<19'b0111010010100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111010010100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0111010010100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111010010100111010) && ({row_reg, col_reg}<19'b0111010010100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111010010100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0111010010100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111010010100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111010010100111111) && ({row_reg, col_reg}<19'b0111010010101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111010010101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0111010010101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0111010010101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0111010010101010100) && ({row_reg, col_reg}<19'b0111010010111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111010010111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0111010010111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111010010111010000) && ({row_reg, col_reg}<19'b0111010010111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111010010111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0111010010111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0111010010111101010) && ({row_reg, col_reg}<19'b0111010100100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111010100100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0111010100100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111010100100111010) && ({row_reg, col_reg}<19'b0111010100100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111010100100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0111010100100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111010100100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111010100100111111) && ({row_reg, col_reg}<19'b0111010100101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111010100101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0111010100101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0111010100101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0111010100101010100) && ({row_reg, col_reg}<19'b0111010100111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111010100111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0111010100111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111010100111010000) && ({row_reg, col_reg}<19'b0111010100111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111010100111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0111010100111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0111010100111101010) && ({row_reg, col_reg}<19'b0111010110100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111010110100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0111010110100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111010110100111010) && ({row_reg, col_reg}<19'b0111010110100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111010110100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0111010110100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111010110100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111010110100111111) && ({row_reg, col_reg}<19'b0111010110101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111010110101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0111010110101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0111010110101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0111010110101010100) && ({row_reg, col_reg}<19'b0111010110111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111010110111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0111010110111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111010110111010000) && ({row_reg, col_reg}<19'b0111010110111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111010110111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0111010110111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0111010110111101010) && ({row_reg, col_reg}<19'b0111011000100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111011000100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0111011000100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111011000100111010) && ({row_reg, col_reg}<19'b0111011000100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111011000100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0111011000100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111011000100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111011000100111111) && ({row_reg, col_reg}<19'b0111011000101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111011000101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0111011000101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0111011000101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0111011000101010100) && ({row_reg, col_reg}<19'b0111011000111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111011000111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0111011000111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111011000111010000) && ({row_reg, col_reg}<19'b0111011000111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111011000111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0111011000111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0111011000111101010) && ({row_reg, col_reg}<19'b0111011010100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111011010100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0111011010100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111011010100111010) && ({row_reg, col_reg}<19'b0111011010100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111011010100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0111011010100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111011010100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111011010100111111) && ({row_reg, col_reg}<19'b0111011010101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111011010101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0111011010101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0111011010101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0111011010101010100) && ({row_reg, col_reg}<19'b0111011010111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111011010111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0111011010111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111011010111010000) && ({row_reg, col_reg}<19'b0111011010111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111011010111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0111011010111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0111011010111101010) && ({row_reg, col_reg}<19'b0111011100100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111011100100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0111011100100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111011100100111010) && ({row_reg, col_reg}<19'b0111011100100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111011100100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0111011100100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111011100100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111011100100111111) && ({row_reg, col_reg}<19'b0111011100101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111011100101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0111011100101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0111011100101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0111011100101010100) && ({row_reg, col_reg}<19'b0111011100111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111011100111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0111011100111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111011100111010000) && ({row_reg, col_reg}<19'b0111011100111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111011100111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0111011100111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0111011100111101010) && ({row_reg, col_reg}<19'b0111011110100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111011110100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0111011110100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111011110100111010) && ({row_reg, col_reg}<19'b0111011110100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111011110100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0111011110100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111011110100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111011110100111111) && ({row_reg, col_reg}<19'b0111011110101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111011110101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0111011110101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0111011110101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0111011110101010100) && ({row_reg, col_reg}<19'b0111011110111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111011110111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0111011110111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111011110111010000) && ({row_reg, col_reg}<19'b0111011110111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111011110111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0111011110111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0111011110111101010) && ({row_reg, col_reg}<19'b0111100000100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111100000100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0111100000100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111100000100111010) && ({row_reg, col_reg}<19'b0111100000100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111100000100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0111100000100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111100000100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111100000100111111) && ({row_reg, col_reg}<19'b0111100000101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111100000101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0111100000101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0111100000101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0111100000101010100) && ({row_reg, col_reg}<19'b0111100000111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111100000111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0111100000111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111100000111010000) && ({row_reg, col_reg}<19'b0111100000111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111100000111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0111100000111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0111100000111101010) && ({row_reg, col_reg}<19'b0111100010100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111100010100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0111100010100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111100010100111010) && ({row_reg, col_reg}<19'b0111100010100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111100010100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0111100010100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111100010100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111100010100111111) && ({row_reg, col_reg}<19'b0111100010101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111100010101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0111100010101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0111100010101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0111100010101010100) && ({row_reg, col_reg}<19'b0111100010111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111100010111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0111100010111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111100010111010000) && ({row_reg, col_reg}<19'b0111100010111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111100010111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0111100010111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0111100010111101010) && ({row_reg, col_reg}<19'b0111100100100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111100100100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0111100100100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111100100100111010) && ({row_reg, col_reg}<19'b0111100100100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111100100100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0111100100100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111100100100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111100100100111111) && ({row_reg, col_reg}<19'b0111100100101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111100100101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0111100100101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0111100100101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0111100100101010100) && ({row_reg, col_reg}<19'b0111100100111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111100100111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0111100100111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111100100111010000) && ({row_reg, col_reg}<19'b0111100100111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111100100111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0111100100111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0111100100111101010) && ({row_reg, col_reg}<19'b0111100110100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111100110100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0111100110100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111100110100111010) && ({row_reg, col_reg}<19'b0111100110100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111100110100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0111100110100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111100110100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111100110100111111) && ({row_reg, col_reg}<19'b0111100110101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111100110101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0111100110101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0111100110101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0111100110101010100) && ({row_reg, col_reg}<19'b0111100110111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111100110111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0111100110111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111100110111010000) && ({row_reg, col_reg}<19'b0111100110111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111100110111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0111100110111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0111100110111101010) && ({row_reg, col_reg}<19'b0111101000100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111101000100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0111101000100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111101000100111010) && ({row_reg, col_reg}<19'b0111101000100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111101000100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0111101000100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111101000100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111101000100111111) && ({row_reg, col_reg}<19'b0111101000101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111101000101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0111101000101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0111101000101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0111101000101010100) && ({row_reg, col_reg}<19'b0111101000111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111101000111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0111101000111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111101000111010000) && ({row_reg, col_reg}<19'b0111101000111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111101000111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0111101000111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0111101000111101010) && ({row_reg, col_reg}<19'b0111101010100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111101010100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0111101010100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111101010100111010) && ({row_reg, col_reg}<19'b0111101010100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111101010100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0111101010100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111101010100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111101010100111111) && ({row_reg, col_reg}<19'b0111101010101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111101010101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0111101010101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0111101010101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0111101010101010100) && ({row_reg, col_reg}<19'b0111101010111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111101010111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0111101010111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111101010111010000) && ({row_reg, col_reg}<19'b0111101010111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111101010111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0111101010111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0111101010111101010) && ({row_reg, col_reg}<19'b0111101100100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111101100100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0111101100100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111101100100111010) && ({row_reg, col_reg}<19'b0111101100100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111101100100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0111101100100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111101100100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111101100100111111) && ({row_reg, col_reg}<19'b0111101100101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111101100101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0111101100101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0111101100101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0111101100101010100) && ({row_reg, col_reg}<19'b0111101100111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111101100111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0111101100111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111101100111010000) && ({row_reg, col_reg}<19'b0111101100111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111101100111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0111101100111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0111101100111101010) && ({row_reg, col_reg}<19'b0111101110100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111101110100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0111101110100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111101110100111010) && ({row_reg, col_reg}<19'b0111101110100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111101110100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0111101110100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111101110100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111101110100111111) && ({row_reg, col_reg}<19'b0111101110101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111101110101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0111101110101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0111101110101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0111101110101010100) && ({row_reg, col_reg}<19'b0111101110111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111101110111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0111101110111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111101110111010000) && ({row_reg, col_reg}<19'b0111101110111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111101110111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0111101110111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0111101110111101010) && ({row_reg, col_reg}<19'b0111110000100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111110000100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0111110000100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111110000100111010) && ({row_reg, col_reg}<19'b0111110000100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111110000100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0111110000100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111110000100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111110000100111111) && ({row_reg, col_reg}<19'b0111110000101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111110000101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0111110000101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0111110000101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0111110000101010100) && ({row_reg, col_reg}<19'b0111110000111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111110000111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0111110000111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111110000111010000) && ({row_reg, col_reg}<19'b0111110000111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111110000111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0111110000111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0111110000111101010) && ({row_reg, col_reg}<19'b0111110010100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111110010100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0111110010100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111110010100111010) && ({row_reg, col_reg}<19'b0111110010100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111110010100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0111110010100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111110010100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111110010100111111) && ({row_reg, col_reg}<19'b0111110010101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111110010101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0111110010101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0111110010101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0111110010101010100) && ({row_reg, col_reg}<19'b0111110010111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111110010111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0111110010111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111110010111010000) && ({row_reg, col_reg}<19'b0111110010111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111110010111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0111110010111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0111110010111101010) && ({row_reg, col_reg}<19'b0111110100100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111110100100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0111110100100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111110100100111010) && ({row_reg, col_reg}<19'b0111110100100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111110100100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0111110100100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111110100100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111110100100111111) && ({row_reg, col_reg}<19'b0111110100101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111110100101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0111110100101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0111110100101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0111110100101010100) && ({row_reg, col_reg}<19'b0111110100111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111110100111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0111110100111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111110100111010000) && ({row_reg, col_reg}<19'b0111110100111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111110100111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0111110100111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0111110100111101010) && ({row_reg, col_reg}<19'b0111110110100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111110110100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0111110110100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111110110100111010) && ({row_reg, col_reg}<19'b0111110110100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111110110100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0111110110100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111110110100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111110110100111111) && ({row_reg, col_reg}<19'b0111110110101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111110110101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0111110110101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0111110110101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0111110110101010100) && ({row_reg, col_reg}<19'b0111110110111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111110110111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0111110110111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111110110111010000) && ({row_reg, col_reg}<19'b0111110110111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111110110111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0111110110111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0111110110111101010) && ({row_reg, col_reg}<19'b0111111000100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111111000100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0111111000100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111111000100111010) && ({row_reg, col_reg}<19'b0111111000100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111111000100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0111111000100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111111000100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111111000100111111) && ({row_reg, col_reg}<19'b0111111000101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111111000101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0111111000101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0111111000101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0111111000101010100) && ({row_reg, col_reg}<19'b0111111000111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111111000111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0111111000111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111111000111010000) && ({row_reg, col_reg}<19'b0111111000111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111111000111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0111111000111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0111111000111101010) && ({row_reg, col_reg}<19'b0111111010100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111111010100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0111111010100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111111010100111010) && ({row_reg, col_reg}<19'b0111111010100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111111010100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0111111010100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111111010100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111111010100111111) && ({row_reg, col_reg}<19'b0111111010101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111111010101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0111111010101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0111111010101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0111111010101010100) && ({row_reg, col_reg}<19'b0111111010111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111111010111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0111111010111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111111010111010000) && ({row_reg, col_reg}<19'b0111111010111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111111010111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0111111010111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0111111010111101010) && ({row_reg, col_reg}<19'b0111111100100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111111100100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0111111100100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111111100100111010) && ({row_reg, col_reg}<19'b0111111100100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111111100100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0111111100100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111111100100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111111100100111111) && ({row_reg, col_reg}<19'b0111111100101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111111100101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0111111100101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0111111100101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0111111100101010100) && ({row_reg, col_reg}<19'b0111111100111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111111100111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0111111100111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111111100111010000) && ({row_reg, col_reg}<19'b0111111100111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111111100111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0111111100111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0111111100111101010) && ({row_reg, col_reg}<19'b0111111110100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111111110100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b0111111110100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111111110100111010) && ({row_reg, col_reg}<19'b0111111110100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111111110100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0111111110100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111111110100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111111110100111111) && ({row_reg, col_reg}<19'b0111111110101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111111110101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b0111111110101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b0111111110101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b0111111110101010100) && ({row_reg, col_reg}<19'b0111111110111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b0111111110111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b0111111110111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b0111111110111010000) && ({row_reg, col_reg}<19'b0111111110111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b0111111110111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b0111111110111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b0111111110111101010) && ({row_reg, col_reg}<19'b1000000000100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000000000100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1000000000100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000000000100111010) && ({row_reg, col_reg}<19'b1000000000100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000000000100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1000000000100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000000000100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000000000100111111) && ({row_reg, col_reg}<19'b1000000000101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000000000101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1000000000101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1000000000101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1000000000101010100) && ({row_reg, col_reg}<19'b1000000000111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000000000111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1000000000111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000000000111010000) && ({row_reg, col_reg}<19'b1000000000111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000000000111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1000000000111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1000000000111101010) && ({row_reg, col_reg}<19'b1000000010100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000000010100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1000000010100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000000010100111010) && ({row_reg, col_reg}<19'b1000000010100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000000010100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1000000010100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000000010100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000000010100111111) && ({row_reg, col_reg}<19'b1000000010101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000000010101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1000000010101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1000000010101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1000000010101010100) && ({row_reg, col_reg}<19'b1000000010111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000000010111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1000000010111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000000010111010000) && ({row_reg, col_reg}<19'b1000000010111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000000010111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1000000010111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1000000010111101010) && ({row_reg, col_reg}<19'b1000000100100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000000100100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1000000100100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000000100100111010) && ({row_reg, col_reg}<19'b1000000100100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000000100100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1000000100100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000000100100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000000100100111111) && ({row_reg, col_reg}<19'b1000000100101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000000100101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1000000100101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1000000100101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1000000100101010100) && ({row_reg, col_reg}<19'b1000000100111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000000100111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1000000100111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000000100111010000) && ({row_reg, col_reg}<19'b1000000100111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000000100111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1000000100111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1000000100111101010) && ({row_reg, col_reg}<19'b1000000110100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000000110100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1000000110100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000000110100111010) && ({row_reg, col_reg}<19'b1000000110100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000000110100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1000000110100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000000110100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000000110100111111) && ({row_reg, col_reg}<19'b1000000110101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000000110101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1000000110101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1000000110101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1000000110101010100) && ({row_reg, col_reg}<19'b1000000110111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000000110111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1000000110111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000000110111010000) && ({row_reg, col_reg}<19'b1000000110111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000000110111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1000000110111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1000000110111101010) && ({row_reg, col_reg}<19'b1000001000100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000001000100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1000001000100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000001000100111010) && ({row_reg, col_reg}<19'b1000001000100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000001000100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1000001000100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000001000100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000001000100111111) && ({row_reg, col_reg}<19'b1000001000101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000001000101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1000001000101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1000001000101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1000001000101010100) && ({row_reg, col_reg}<19'b1000001000111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000001000111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1000001000111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000001000111010000) && ({row_reg, col_reg}<19'b1000001000111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000001000111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1000001000111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1000001000111101010) && ({row_reg, col_reg}<19'b1000001010100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000001010100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1000001010100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000001010100111010) && ({row_reg, col_reg}<19'b1000001010100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000001010100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1000001010100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000001010100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000001010100111111) && ({row_reg, col_reg}<19'b1000001010101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000001010101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1000001010101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1000001010101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1000001010101010100) && ({row_reg, col_reg}<19'b1000001010111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000001010111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1000001010111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000001010111010000) && ({row_reg, col_reg}<19'b1000001010111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000001010111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1000001010111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1000001010111101010) && ({row_reg, col_reg}<19'b1000001100100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000001100100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1000001100100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000001100100111010) && ({row_reg, col_reg}<19'b1000001100100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000001100100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1000001100100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000001100100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000001100100111111) && ({row_reg, col_reg}<19'b1000001100101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000001100101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1000001100101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1000001100101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1000001100101010100) && ({row_reg, col_reg}<19'b1000001100111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000001100111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1000001100111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000001100111010000) && ({row_reg, col_reg}<19'b1000001100111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000001100111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1000001100111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1000001100111101010) && ({row_reg, col_reg}<19'b1000001110100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000001110100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1000001110100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000001110100111010) && ({row_reg, col_reg}<19'b1000001110100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000001110100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1000001110100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000001110100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000001110100111111) && ({row_reg, col_reg}<19'b1000001110101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000001110101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1000001110101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1000001110101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1000001110101010100) && ({row_reg, col_reg}<19'b1000001110111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000001110111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1000001110111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000001110111010000) && ({row_reg, col_reg}<19'b1000001110111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000001110111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1000001110111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1000001110111101010) && ({row_reg, col_reg}<19'b1000010000100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000010000100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1000010000100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000010000100111010) && ({row_reg, col_reg}<19'b1000010000100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000010000100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1000010000100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000010000100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000010000100111111) && ({row_reg, col_reg}<19'b1000010000101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000010000101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1000010000101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1000010000101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1000010000101010100) && ({row_reg, col_reg}<19'b1000010000111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000010000111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1000010000111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000010000111010000) && ({row_reg, col_reg}<19'b1000010000111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000010000111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1000010000111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1000010000111101010) && ({row_reg, col_reg}<19'b1000010010100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000010010100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1000010010100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000010010100111010) && ({row_reg, col_reg}<19'b1000010010100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000010010100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1000010010100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000010010100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000010010100111111) && ({row_reg, col_reg}<19'b1000010010101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000010010101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1000010010101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1000010010101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1000010010101010100) && ({row_reg, col_reg}<19'b1000010010111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000010010111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1000010010111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000010010111010000) && ({row_reg, col_reg}<19'b1000010010111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000010010111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1000010010111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1000010010111101010) && ({row_reg, col_reg}<19'b1000010100100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000010100100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1000010100100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000010100100111010) && ({row_reg, col_reg}<19'b1000010100100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000010100100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1000010100100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000010100100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000010100100111111) && ({row_reg, col_reg}<19'b1000010100101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000010100101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1000010100101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1000010100101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1000010100101010100) && ({row_reg, col_reg}<19'b1000010100111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000010100111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1000010100111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000010100111010000) && ({row_reg, col_reg}<19'b1000010100111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000010100111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1000010100111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1000010100111101010) && ({row_reg, col_reg}<19'b1000010110100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000010110100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1000010110100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000010110100111010) && ({row_reg, col_reg}<19'b1000010110100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000010110100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1000010110100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000010110100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000010110100111111) && ({row_reg, col_reg}<19'b1000010110101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000010110101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1000010110101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1000010110101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1000010110101010100) && ({row_reg, col_reg}<19'b1000010110111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000010110111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1000010110111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000010110111010000) && ({row_reg, col_reg}<19'b1000010110111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000010110111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1000010110111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1000010110111101010) && ({row_reg, col_reg}<19'b1000011000100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000011000100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1000011000100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000011000100111010) && ({row_reg, col_reg}<19'b1000011000100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000011000100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1000011000100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000011000100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000011000100111111) && ({row_reg, col_reg}<19'b1000011000101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000011000101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1000011000101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1000011000101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1000011000101010100) && ({row_reg, col_reg}<19'b1000011000111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000011000111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1000011000111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000011000111010000) && ({row_reg, col_reg}<19'b1000011000111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000011000111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1000011000111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1000011000111101010) && ({row_reg, col_reg}<19'b1000011010100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000011010100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1000011010100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000011010100111010) && ({row_reg, col_reg}<19'b1000011010100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000011010100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1000011010100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000011010100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000011010100111111) && ({row_reg, col_reg}<19'b1000011010101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000011010101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1000011010101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1000011010101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1000011010101010100) && ({row_reg, col_reg}<19'b1000011010111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000011010111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1000011010111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000011010111010000) && ({row_reg, col_reg}<19'b1000011010111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000011010111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1000011010111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1000011010111101010) && ({row_reg, col_reg}<19'b1000011100100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000011100100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1000011100100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000011100100111010) && ({row_reg, col_reg}<19'b1000011100100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000011100100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1000011100100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000011100100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000011100100111111) && ({row_reg, col_reg}<19'b1000011100101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000011100101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1000011100101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1000011100101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1000011100101010100) && ({row_reg, col_reg}<19'b1000011100111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000011100111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1000011100111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000011100111010000) && ({row_reg, col_reg}<19'b1000011100111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000011100111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1000011100111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1000011100111101010) && ({row_reg, col_reg}<19'b1000011110100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000011110100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1000011110100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000011110100111010) && ({row_reg, col_reg}<19'b1000011110100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000011110100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1000011110100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000011110100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000011110100111111) && ({row_reg, col_reg}<19'b1000011110101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000011110101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1000011110101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1000011110101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1000011110101010100) && ({row_reg, col_reg}<19'b1000011110111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000011110111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1000011110111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000011110111010000) && ({row_reg, col_reg}<19'b1000011110111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000011110111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1000011110111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1000011110111101010) && ({row_reg, col_reg}<19'b1000100000100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000100000100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1000100000100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000100000100111010) && ({row_reg, col_reg}<19'b1000100000100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000100000100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1000100000100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000100000100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000100000100111111) && ({row_reg, col_reg}<19'b1000100000101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000100000101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1000100000101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1000100000101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1000100000101010100) && ({row_reg, col_reg}<19'b1000100000111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000100000111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1000100000111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000100000111010000) && ({row_reg, col_reg}<19'b1000100000111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000100000111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1000100000111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1000100000111101010) && ({row_reg, col_reg}<19'b1000100010100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000100010100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1000100010100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000100010100111010) && ({row_reg, col_reg}<19'b1000100010100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000100010100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1000100010100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000100010100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000100010100111111) && ({row_reg, col_reg}<19'b1000100010101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000100010101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1000100010101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1000100010101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1000100010101010100) && ({row_reg, col_reg}<19'b1000100010111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000100010111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1000100010111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000100010111010000) && ({row_reg, col_reg}<19'b1000100010111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000100010111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1000100010111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1000100010111101010) && ({row_reg, col_reg}<19'b1000100100100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000100100100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1000100100100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000100100100111010) && ({row_reg, col_reg}<19'b1000100100100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000100100100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1000100100100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000100100100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000100100100111111) && ({row_reg, col_reg}<19'b1000100100101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000100100101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1000100100101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1000100100101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1000100100101010100) && ({row_reg, col_reg}<19'b1000100100111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000100100111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1000100100111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000100100111010000) && ({row_reg, col_reg}<19'b1000100100111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000100100111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1000100100111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1000100100111101010) && ({row_reg, col_reg}<19'b1000100110100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000100110100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1000100110100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000100110100111010) && ({row_reg, col_reg}<19'b1000100110100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000100110100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1000100110100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000100110100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000100110100111111) && ({row_reg, col_reg}<19'b1000100110101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000100110101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1000100110101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1000100110101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1000100110101010100) && ({row_reg, col_reg}<19'b1000100110111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000100110111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1000100110111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000100110111010000) && ({row_reg, col_reg}<19'b1000100110111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000100110111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1000100110111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1000100110111101010) && ({row_reg, col_reg}<19'b1000101000100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000101000100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1000101000100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000101000100111010) && ({row_reg, col_reg}<19'b1000101000100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000101000100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1000101000100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000101000100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000101000100111111) && ({row_reg, col_reg}<19'b1000101000101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000101000101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1000101000101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1000101000101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1000101000101010100) && ({row_reg, col_reg}<19'b1000101000111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000101000111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1000101000111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000101000111010000) && ({row_reg, col_reg}<19'b1000101000111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000101000111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1000101000111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1000101000111101010) && ({row_reg, col_reg}<19'b1000101010100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000101010100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1000101010100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000101010100111010) && ({row_reg, col_reg}<19'b1000101010100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000101010100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1000101010100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000101010100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000101010100111111) && ({row_reg, col_reg}<19'b1000101010101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000101010101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1000101010101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1000101010101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1000101010101010100) && ({row_reg, col_reg}<19'b1000101010111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000101010111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1000101010111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000101010111010000) && ({row_reg, col_reg}<19'b1000101010111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000101010111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1000101010111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1000101010111101010) && ({row_reg, col_reg}<19'b1000101100100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000101100100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1000101100100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000101100100111010) && ({row_reg, col_reg}<19'b1000101100100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000101100100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1000101100100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000101100100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000101100100111111) && ({row_reg, col_reg}<19'b1000101100101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000101100101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1000101100101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1000101100101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1000101100101010100) && ({row_reg, col_reg}<19'b1000101100111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000101100111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1000101100111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000101100111010000) && ({row_reg, col_reg}<19'b1000101100111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000101100111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1000101100111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1000101100111101010) && ({row_reg, col_reg}<19'b1000101110100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000101110100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1000101110100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000101110100111010) && ({row_reg, col_reg}<19'b1000101110100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000101110100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1000101110100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000101110100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000101110100111111) && ({row_reg, col_reg}<19'b1000101110101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000101110101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1000101110101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1000101110101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1000101110101010100) && ({row_reg, col_reg}<19'b1000101110111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000101110111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1000101110111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000101110111010000) && ({row_reg, col_reg}<19'b1000101110111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000101110111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1000101110111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1000101110111101010) && ({row_reg, col_reg}<19'b1000110000100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000110000100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1000110000100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000110000100111010) && ({row_reg, col_reg}<19'b1000110000100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000110000100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1000110000100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000110000100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000110000100111111) && ({row_reg, col_reg}<19'b1000110000101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000110000101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1000110000101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1000110000101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1000110000101010100) && ({row_reg, col_reg}<19'b1000110000111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000110000111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1000110000111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000110000111010000) && ({row_reg, col_reg}<19'b1000110000111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000110000111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1000110000111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1000110000111101010) && ({row_reg, col_reg}<19'b1000110010100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000110010100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1000110010100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000110010100111010) && ({row_reg, col_reg}<19'b1000110010100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000110010100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1000110010100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000110010100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000110010100111111) && ({row_reg, col_reg}<19'b1000110010101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000110010101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1000110010101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1000110010101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1000110010101010100) && ({row_reg, col_reg}<19'b1000110010111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000110010111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1000110010111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000110010111010000) && ({row_reg, col_reg}<19'b1000110010111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000110010111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1000110010111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1000110010111101010) && ({row_reg, col_reg}<19'b1000110100100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000110100100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1000110100100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000110100100111010) && ({row_reg, col_reg}<19'b1000110100100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000110100100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1000110100100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000110100100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000110100100111111) && ({row_reg, col_reg}<19'b1000110100101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000110100101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1000110100101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1000110100101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1000110100101010100) && ({row_reg, col_reg}<19'b1000110100111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000110100111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1000110100111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000110100111010000) && ({row_reg, col_reg}<19'b1000110100111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000110100111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1000110100111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1000110100111101010) && ({row_reg, col_reg}<19'b1000110110100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000110110100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1000110110100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000110110100111010) && ({row_reg, col_reg}<19'b1000110110100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000110110100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1000110110100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000110110100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000110110100111111) && ({row_reg, col_reg}<19'b1000110110101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000110110101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1000110110101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1000110110101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1000110110101010100) && ({row_reg, col_reg}<19'b1000110110111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000110110111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1000110110111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000110110111010000) && ({row_reg, col_reg}<19'b1000110110111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000110110111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1000110110111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1000110110111101010) && ({row_reg, col_reg}<19'b1000111000100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000111000100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1000111000100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000111000100111010) && ({row_reg, col_reg}<19'b1000111000100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000111000100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1000111000100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000111000100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000111000100111111) && ({row_reg, col_reg}<19'b1000111000101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000111000101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1000111000101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1000111000101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1000111000101010100) && ({row_reg, col_reg}<19'b1000111000111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000111000111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1000111000111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000111000111010000) && ({row_reg, col_reg}<19'b1000111000111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000111000111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1000111000111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1000111000111101010) && ({row_reg, col_reg}<19'b1000111010100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000111010100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1000111010100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000111010100111010) && ({row_reg, col_reg}<19'b1000111010100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000111010100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1000111010100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000111010100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000111010100111111) && ({row_reg, col_reg}<19'b1000111010101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000111010101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1000111010101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1000111010101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1000111010101010100) && ({row_reg, col_reg}<19'b1000111010111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000111010111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1000111010111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000111010111010000) && ({row_reg, col_reg}<19'b1000111010111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000111010111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1000111010111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1000111010111101010) && ({row_reg, col_reg}<19'b1000111100100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000111100100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1000111100100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000111100100111010) && ({row_reg, col_reg}<19'b1000111100100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000111100100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1000111100100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000111100100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000111100100111111) && ({row_reg, col_reg}<19'b1000111100101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000111100101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1000111100101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1000111100101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1000111100101010100) && ({row_reg, col_reg}<19'b1000111100111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000111100111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1000111100111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000111100111010000) && ({row_reg, col_reg}<19'b1000111100111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000111100111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1000111100111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1000111100111101010) && ({row_reg, col_reg}<19'b1000111110100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000111110100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1000111110100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000111110100111010) && ({row_reg, col_reg}<19'b1000111110100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000111110100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1000111110100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000111110100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000111110100111111) && ({row_reg, col_reg}<19'b1000111110101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000111110101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1000111110101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1000111110101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1000111110101010100) && ({row_reg, col_reg}<19'b1000111110111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1000111110111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1000111110111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1000111110111010000) && ({row_reg, col_reg}<19'b1000111110111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1000111110111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1000111110111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1000111110111101010) && ({row_reg, col_reg}<19'b1001000000100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1001000000100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1001000000100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001000000100111010) && ({row_reg, col_reg}<19'b1001000000100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001000000100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1001000000100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001000000100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001000000100111111) && ({row_reg, col_reg}<19'b1001000000101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001000000101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1001000000101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1001000000101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1001000000101010100) && ({row_reg, col_reg}<19'b1001000000111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1001000000111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1001000000111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001000000111010000) && ({row_reg, col_reg}<19'b1001000000111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001000000111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1001000000111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1001000000111101010) && ({row_reg, col_reg}<19'b1001000010100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1001000010100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1001000010100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001000010100111010) && ({row_reg, col_reg}<19'b1001000010100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001000010100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1001000010100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001000010100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001000010100111111) && ({row_reg, col_reg}<19'b1001000010101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001000010101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1001000010101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1001000010101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1001000010101010100) && ({row_reg, col_reg}<19'b1001000010111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1001000010111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1001000010111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001000010111010000) && ({row_reg, col_reg}<19'b1001000010111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001000010111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1001000010111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1001000010111101010) && ({row_reg, col_reg}<19'b1001000100100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1001000100100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1001000100100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001000100100111010) && ({row_reg, col_reg}<19'b1001000100100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001000100100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1001000100100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001000100100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001000100100111111) && ({row_reg, col_reg}<19'b1001000100101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001000100101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1001000100101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1001000100101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1001000100101010100) && ({row_reg, col_reg}<19'b1001000100111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1001000100111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1001000100111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001000100111010000) && ({row_reg, col_reg}<19'b1001000100111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001000100111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1001000100111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1001000100111101010) && ({row_reg, col_reg}<19'b1001000110100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1001000110100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1001000110100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001000110100111010) && ({row_reg, col_reg}<19'b1001000110100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001000110100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1001000110100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001000110100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001000110100111111) && ({row_reg, col_reg}<19'b1001000110101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001000110101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1001000110101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1001000110101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1001000110101010100) && ({row_reg, col_reg}<19'b1001000110111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1001000110111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1001000110111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001000110111010000) && ({row_reg, col_reg}<19'b1001000110111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001000110111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1001000110111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1001000110111101010) && ({row_reg, col_reg}<19'b1001001000100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1001001000100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1001001000100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001001000100111010) && ({row_reg, col_reg}<19'b1001001000100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001001000100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1001001000100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001001000100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001001000100111111) && ({row_reg, col_reg}<19'b1001001000101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001001000101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1001001000101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1001001000101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1001001000101010100) && ({row_reg, col_reg}<19'b1001001000111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1001001000111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1001001000111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001001000111010000) && ({row_reg, col_reg}<19'b1001001000111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001001000111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1001001000111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1001001000111101010) && ({row_reg, col_reg}<19'b1001001010100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1001001010100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1001001010100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001001010100111010) && ({row_reg, col_reg}<19'b1001001010100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001001010100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1001001010100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001001010100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001001010100111111) && ({row_reg, col_reg}<19'b1001001010101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001001010101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1001001010101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1001001010101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1001001010101010100) && ({row_reg, col_reg}<19'b1001001010111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1001001010111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1001001010111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001001010111010000) && ({row_reg, col_reg}<19'b1001001010111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001001010111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1001001010111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1001001010111101010) && ({row_reg, col_reg}<19'b1001001100100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1001001100100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1001001100100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001001100100111010) && ({row_reg, col_reg}<19'b1001001100100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001001100100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1001001100100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001001100100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001001100100111111) && ({row_reg, col_reg}<19'b1001001100101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001001100101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1001001100101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1001001100101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1001001100101010100) && ({row_reg, col_reg}<19'b1001001100111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1001001100111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1001001100111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001001100111010000) && ({row_reg, col_reg}<19'b1001001100111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001001100111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1001001100111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1001001100111101010) && ({row_reg, col_reg}<19'b1001001110100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1001001110100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1001001110100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001001110100111010) && ({row_reg, col_reg}<19'b1001001110100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001001110100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1001001110100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001001110100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001001110100111111) && ({row_reg, col_reg}<19'b1001001110101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001001110101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1001001110101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1001001110101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1001001110101010100) && ({row_reg, col_reg}<19'b1001001110111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1001001110111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1001001110111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001001110111010000) && ({row_reg, col_reg}<19'b1001001110111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001001110111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1001001110111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1001001110111101010) && ({row_reg, col_reg}<19'b1001010000100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1001010000100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1001010000100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001010000100111010) && ({row_reg, col_reg}<19'b1001010000100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001010000100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1001010000100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001010000100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001010000100111111) && ({row_reg, col_reg}<19'b1001010000101010000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001010000101010000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1001010000101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001010000101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1001010000101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1001010000101010100) && ({row_reg, col_reg}<19'b1001010000111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1001010000111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1001010000111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001010000111010000) && ({row_reg, col_reg}<19'b1001010000111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001010000111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1001010000111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1001010000111101010) && ({row_reg, col_reg}<19'b1001010010100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1001010010100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1001010010100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001010010100111010) && ({row_reg, col_reg}<19'b1001010010100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001010010100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1001010010100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001010010100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001010010100111111) && ({row_reg, col_reg}<19'b1001010010101010000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001010010101010000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1001010010101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001010010101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1001010010101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1001010010101010100) && ({row_reg, col_reg}<19'b1001010010111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1001010010111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1001010010111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001010010111010000) && ({row_reg, col_reg}<19'b1001010010111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001010010111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1001010010111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1001010010111101010) && ({row_reg, col_reg}<19'b1001010100100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1001010100100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1001010100100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001010100100111010) && ({row_reg, col_reg}<19'b1001010100100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001010100100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1001010100100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001010100100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001010100100111111) && ({row_reg, col_reg}<19'b1001010100101010000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001010100101010000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1001010100101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001010100101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1001010100101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1001010100101010100) && ({row_reg, col_reg}<19'b1001010100111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1001010100111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1001010100111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001010100111010000) && ({row_reg, col_reg}<19'b1001010100111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001010100111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1001010100111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1001010100111101010) && ({row_reg, col_reg}<19'b1001010110100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1001010110100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1001010110100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001010110100111010) && ({row_reg, col_reg}<19'b1001010110100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001010110100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1001010110100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001010110100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001010110100111111) && ({row_reg, col_reg}<19'b1001010110101010000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001010110101010000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1001010110101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001010110101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1001010110101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1001010110101010100) && ({row_reg, col_reg}<19'b1001010110111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1001010110111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1001010110111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001010110111010000) && ({row_reg, col_reg}<19'b1001010110111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001010110111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1001010110111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1001010110111101010) && ({row_reg, col_reg}<19'b1001011000100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1001011000100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1001011000100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001011000100111010) && ({row_reg, col_reg}<19'b1001011000100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001011000100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1001011000100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001011000100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001011000100111111) && ({row_reg, col_reg}<19'b1001011000101010000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001011000101010000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1001011000101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001011000101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1001011000101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1001011000101010100) && ({row_reg, col_reg}<19'b1001011000111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1001011000111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1001011000111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001011000111010000) && ({row_reg, col_reg}<19'b1001011000111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001011000111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1001011000111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1001011000111101010) && ({row_reg, col_reg}<19'b1001011010100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1001011010100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1001011010100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001011010100111010) && ({row_reg, col_reg}<19'b1001011010100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001011010100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1001011010100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001011010100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001011010100111111) && ({row_reg, col_reg}<19'b1001011010101010000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001011010101010000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1001011010101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001011010101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1001011010101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1001011010101010100) && ({row_reg, col_reg}<19'b1001011010111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1001011010111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1001011010111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001011010111010000) && ({row_reg, col_reg}<19'b1001011010111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001011010111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1001011010111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1001011010111101010) && ({row_reg, col_reg}<19'b1001011100100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1001011100100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1001011100100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001011100100111010) && ({row_reg, col_reg}<19'b1001011100100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001011100100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1001011100100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001011100100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001011100100111111) && ({row_reg, col_reg}<19'b1001011100101010000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001011100101010000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1001011100101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001011100101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1001011100101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1001011100101010100) && ({row_reg, col_reg}<19'b1001011100111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1001011100111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1001011100111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001011100111010000) && ({row_reg, col_reg}<19'b1001011100111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001011100111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1001011100111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1001011100111101010) && ({row_reg, col_reg}<19'b1001011110100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1001011110100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1001011110100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001011110100111010) && ({row_reg, col_reg}<19'b1001011110100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001011110100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1001011110100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001011110100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001011110100111111) && ({row_reg, col_reg}<19'b1001011110101010000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001011110101010000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1001011110101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001011110101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1001011110101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1001011110101010100) && ({row_reg, col_reg}<19'b1001011110111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1001011110111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1001011110111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001011110111010000) && ({row_reg, col_reg}<19'b1001011110111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001011110111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1001011110111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1001011110111101010) && ({row_reg, col_reg}<19'b1001100000100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1001100000100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1001100000100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1001100000100111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001100000100111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001100000100111100) && ({row_reg, col_reg}<19'b1001100000101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001100000101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1001100000101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1001100000101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1001100000101010100) && ({row_reg, col_reg}<19'b1001100000111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1001100000111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1001100000111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001100000111010000) && ({row_reg, col_reg}<19'b1001100000111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001100000111101000)) color_data = 12'b101010101010;

		if(({row_reg, col_reg}>=19'b1001100000111101001) && ({row_reg, col_reg}<19'b1001100010100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1001100010100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1001100010100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001100010100111010) && ({row_reg, col_reg}<19'b1001100010101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001100010101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1001100010101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1001100010101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1001100010101010100) && ({row_reg, col_reg}<19'b1001100010111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1001100010111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1001100010111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001100010111010000) && ({row_reg, col_reg}<19'b1001100010111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001100010111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1001100010111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1001100010111101010) && ({row_reg, col_reg}<19'b1001100100010101001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1001100100010101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=19'b1001100100010101010) && ({row_reg, col_reg}<19'b1001100100010101100)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1001100100010101100) && ({row_reg, col_reg}<19'b1001100100010101110)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=19'b1001100100010101110) && ({row_reg, col_reg}<19'b1001100100100111000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1001100100100111000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1001100100100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001100100100111010) && ({row_reg, col_reg}<19'b1001100100100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001100100100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1001100100100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001100100100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001100100100111111) && ({row_reg, col_reg}<19'b1001100100101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b1001100100101010001) && ({row_reg, col_reg}<19'b1001100100101010011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1001100100101010011)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=19'b1001100100101010100) && ({row_reg, col_reg}<19'b1001100100111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1001100100111001110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=19'b1001100100111001111) && ({row_reg, col_reg}<19'b1001100100111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001100100111101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001100100111101001) && ({row_reg, col_reg}<19'b1001100101001110001)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=19'b1001100101001110001) && ({row_reg, col_reg}<19'b1001100101001110011)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1001100101001110011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1001100101001110100) && ({row_reg, col_reg}<19'b1001100101001110110)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1001100101001110110) && ({row_reg, col_reg}<19'b1001100110010100110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1001100110010100110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b1001100110010100111)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b1001100110010101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1001100110010101001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1001100110010101010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=19'b1001100110010101011) && ({row_reg, col_reg}<19'b1001100110010101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1001100110010101110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b1001100110010101111) && ({row_reg, col_reg}<19'b1001100110100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001100110100111001) && ({row_reg, col_reg}<19'b1001100110100111011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b1001100110100111011) && ({row_reg, col_reg}<19'b1001100110100111101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1001100110100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001100110100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001100110100111111) && ({row_reg, col_reg}<19'b1001100110101010000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b1001100110101010000) && ({row_reg, col_reg}<19'b1001100110101010010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1001100110101010010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b1001100110101010011) && ({row_reg, col_reg}<19'b1001100110111010000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001100110111010000) && ({row_reg, col_reg}<19'b1001100110111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b1001100110111101000) && ({row_reg, col_reg}<19'b1001100111001110011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001100111001110011) && ({row_reg, col_reg}<19'b1001100111001110101)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1001100111001110101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1001100111001110110)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1001100111001110111)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1001100111001111000) && ({row_reg, col_reg}<19'b1001101000010100101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1001101000010100101)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b1001101000010100110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1001101000010100111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1001101000010101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001101000010101001) && ({row_reg, col_reg}<19'b1001101000010101011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b1001101000010101011) && ({row_reg, col_reg}<19'b1001101000010110000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001101000010110000) && ({row_reg, col_reg}<19'b1001101000100111001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001101000100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1001101000100111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001101000100111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001101000100111100) && ({row_reg, col_reg}<19'b1001101000100111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b1001101000100111110) && ({row_reg, col_reg}<19'b1001101000101000000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001101000101000000) && ({row_reg, col_reg}<19'b1001101000101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001101000101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1001101000101010010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001101000101010011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1001101000101010100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001101000101010101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001101000101010110) && ({row_reg, col_reg}<19'b1001101000111001000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b1001101000111001000) && ({row_reg, col_reg}<19'b1001101000111001010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001101000111001010) && ({row_reg, col_reg}<19'b1001101000111001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001101000111001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001101000111001101) && ({row_reg, col_reg}<19'b1001101000111101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001101000111101101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001101000111101110) && ({row_reg, col_reg}<19'b1001101001001110000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001101001001110000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001101001001110001) && ({row_reg, col_reg}<19'b1001101001001110110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001101001001110110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1001101001001110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1001101001001111000)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b1001101001001111001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1001101001001111010) && ({row_reg, col_reg}<19'b1001101010010100100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1001101010010100100)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b1001101010010100101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1001101010010100110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001101010010100111) && ({row_reg, col_reg}<19'b1001101010010101011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b1001101010010101011) && ({row_reg, col_reg}<19'b1001101010010101101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001101010010101101) && ({row_reg, col_reg}<19'b1001101010010110000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b1001101010010110000) && ({row_reg, col_reg}<19'b1001101010100111000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1001101010100111000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001101010100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1001101010100111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001101010100111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1001101010100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001101010100111101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001101010100111110) && ({row_reg, col_reg}<19'b1001101010101010010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001101010101010010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001101010101010011) && ({row_reg, col_reg}<19'b1001101010101011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b1001101010101011000) && ({row_reg, col_reg}<19'b1001101010111001001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001101010111001001) && ({row_reg, col_reg}<19'b1001101010111001011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b1001101010111001011) && ({row_reg, col_reg}<19'b1001101010111001101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001101010111001101) && ({row_reg, col_reg}<19'b1001101010111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b1001101010111101000) && ({row_reg, col_reg}<19'b1001101010111101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1001101010111101110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b1001101010111101111) && ({row_reg, col_reg}<19'b1001101011001110000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001101011001110000) && ({row_reg, col_reg}<19'b1001101011001110111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001101011001110111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1001101011001111000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1001101011001111001)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1001101011001111010)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1001101011001111011) && ({row_reg, col_reg}<19'b1001101100010100011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1001101100010100011)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1001101100010100100)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=19'b1001101100010100101) && ({row_reg, col_reg}<19'b1001101100010100111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b1001101100010100111) && ({row_reg, col_reg}<19'b1001101100010101011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001101100010101011) && ({row_reg, col_reg}<19'b1001101100010101110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b1001101100010101110) && ({row_reg, col_reg}<19'b1001101100010110000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001101100010110000) && ({row_reg, col_reg}<19'b1001101100100111011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001101100100111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1001101100100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001101100100111101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001101100100111110) && ({row_reg, col_reg}<19'b1001101100101010000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b1001101100101010000) && ({row_reg, col_reg}<19'b1001101100101010011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001101100101010011) && ({row_reg, col_reg}<19'b1001101100101010101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b1001101100101010101) && ({row_reg, col_reg}<19'b1001101100101011000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001101100101011000) && ({row_reg, col_reg}<19'b1001101100111001011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001101100111001011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1001101100111001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b1001101100111001101) && ({row_reg, col_reg}<19'b1001101100111010000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001101100111010000) && ({row_reg, col_reg}<19'b1001101100111101110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b1001101100111101110) && ({row_reg, col_reg}<19'b1001101100111110000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001101100111110000) && ({row_reg, col_reg}<19'b1001101101001110000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b1001101101001110000) && ({row_reg, col_reg}<19'b1001101101001110011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001101101001110011) && ({row_reg, col_reg}<19'b1001101101001110101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b1001101101001110101) && ({row_reg, col_reg}<19'b1001101101001110111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001101101001110111) && ({row_reg, col_reg}<19'b1001101101001111001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001101101001111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1001101101001111010)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1001101101001111011)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1001101101001111100) && ({row_reg, col_reg}<19'b1001101110010100010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1001101110010100010)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b1001101110010100011)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=19'b1001101110010100100) && ({row_reg, col_reg}<19'b1001101110010100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001101110010100110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001101110010100111) && ({row_reg, col_reg}<19'b1001101110010101010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001101110010101010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001101110010101011) && ({row_reg, col_reg}<19'b1001101110010101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b1001101110010101101) && ({row_reg, col_reg}<19'b1001101110010101111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001101110010101111) && ({row_reg, col_reg}<19'b1001101110100111011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001101110100111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1001101110100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001101110100111101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1001101110100111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001101110100111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001101110101000000) && ({row_reg, col_reg}<19'b1001101110101010000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001101110101010000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001101110101010001) && ({row_reg, col_reg}<19'b1001101110101010100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b1001101110101010100) && ({row_reg, col_reg}<19'b1001101110101010110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001101110101010110) && ({row_reg, col_reg}<19'b1001101110111001000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b1001101110111001000) && ({row_reg, col_reg}<19'b1001101110111001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1001101110111001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001101110111001101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001101110111001110) && ({row_reg, col_reg}<19'b1001101110111101001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001101110111101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001101110111101010) && ({row_reg, col_reg}<19'b1001101110111101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b1001101110111101100) && ({row_reg, col_reg}<19'b1001101110111101111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001101110111101111) && ({row_reg, col_reg}<19'b1001101111001111000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001101111001111000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1001101111001111001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001101111001111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1001101111001111011)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=19'b1001101111001111100) && ({row_reg, col_reg}<19'b1001110000010100001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1001110000010100001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b1001110000010100010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1001110000010100011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001110000010100100) && ({row_reg, col_reg}<19'b1001110000010100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001110000010100110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001110000010100111) && ({row_reg, col_reg}<19'b1001110001001111001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b1001110001001111001) && ({row_reg, col_reg}<19'b1001110001001111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1001110001001111100)) color_data = 12'b110111011101;

		if(({row_reg, col_reg}>=19'b1001110001001111101) && ({row_reg, col_reg}<19'b1001110010010100001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1001110010010100001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1001110010010100010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1001110010010100011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001110010010100100) && ({row_reg, col_reg}<19'b1001110010010100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001110010010100110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001110010010100111) && ({row_reg, col_reg}<19'b1001110011001111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001110011001111100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1001110011001111101)) color_data = 12'b110111011101;

		if(({row_reg, col_reg}>=19'b1001110011001111110) && ({row_reg, col_reg}<19'b1001110100010100000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1001110100010100000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b1001110100010100001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=19'b1001110100010100010) && ({row_reg, col_reg}<19'b1001110100010100100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b1001110100010100100) && ({row_reg, col_reg}<19'b1001110100010100111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001110100010100111) && ({row_reg, col_reg}<19'b1001110101001111000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001110101001111000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001110101001111001) && ({row_reg, col_reg}<19'b1001110101001111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001110101001111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1001110101001111101)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=19'b1001110101001111110) && ({row_reg, col_reg}<19'b1001110110010100000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1001110110010100000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1001110110010100001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1001110110010100010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001110110010100011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1001110110010100100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b1001110110010100101) && ({row_reg, col_reg}<19'b1001110110010100111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001110110010100111) && ({row_reg, col_reg}<19'b1001110111001111001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b1001110111001111001) && ({row_reg, col_reg}<19'b1001110111001111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1001110111001111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001110111001111101)) color_data = 12'b101110111011;

		if(({row_reg, col_reg}>=19'b1001110111001111110) && ({row_reg, col_reg}<19'b1001111000010100000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1001111000010100000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1001111000010100001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1001111000010100010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001111000010100011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1001111000010100100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001111000010100101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001111000010100110) && ({row_reg, col_reg}<19'b1001111001001111001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b1001111001001111001) && ({row_reg, col_reg}<19'b1001111001001111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1001111001001111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001111001001111101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1001111001001111110)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1001111001001111111) && ({row_reg, col_reg}<19'b1001111010010100000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1001111010010100000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1001111010010100001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1001111010010100010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001111010010100011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001111010010100100) && ({row_reg, col_reg}<19'b1001111010010100111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001111010010100111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001111010010101000) && ({row_reg, col_reg}<19'b1001111011001111000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b1001111011001111000) && ({row_reg, col_reg}<19'b1001111011001111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001111011001111010) && ({row_reg, col_reg}<19'b1001111011001111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001111011001111101)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1001111011001111110)) color_data = 12'b110111011101;

		if(({row_reg, col_reg}>=19'b1001111011001111111) && ({row_reg, col_reg}<19'b1001111100010100000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1001111100010100000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1001111100010100001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001111100010100010) && ({row_reg, col_reg}<19'b1001111100010100100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b1001111100010100100) && ({row_reg, col_reg}<19'b1001111100010100110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1001111100010100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001111100010100111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001111100010101000) && ({row_reg, col_reg}<19'b1001111101001111000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001111101001111000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1001111101001111001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001111101001111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001111101001111011) && ({row_reg, col_reg}<19'b1001111101001111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001111101001111101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1001111101001111110)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=19'b1001111101001111111) && ({row_reg, col_reg}<19'b1001111110010100000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=19'b1001111110010100000) && ({row_reg, col_reg}<19'b1001111110010100010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001111110010100010) && ({row_reg, col_reg}<19'b1001111110010100100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b1001111110010100100) && ({row_reg, col_reg}<19'b1001111110010100110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001111110010100110) && ({row_reg, col_reg}<19'b1001111111001111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001111111001111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1001111111001111011) && ({row_reg, col_reg}<19'b1001111111001111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1001111111001111101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1001111111001111110)) color_data = 12'b101110111011;

		if(({row_reg, col_reg}>=19'b1001111111001111111) && ({row_reg, col_reg}<19'b1010000000010100000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=19'b1010000000010100000) && ({row_reg, col_reg}<19'b1010000000010100010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1010000000010100010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010000000010100011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1010000000010100100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b1010000000010100101) && ({row_reg, col_reg}<19'b1010000000010100111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010000000010100111) && ({row_reg, col_reg}<19'b1010000001001111000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010000001001111000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1010000001001111001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010000001001111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010000001001111011) && ({row_reg, col_reg}<19'b1010000001001111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010000001001111101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1010000001001111110)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=19'b1010000001001111111) && ({row_reg, col_reg}<19'b1010000010010100000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1010000010010100000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1010000010010100001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010000010010100010) && ({row_reg, col_reg}<19'b1010000010010100101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b1010000010010100101) && ({row_reg, col_reg}<19'b1010000010010101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010000010010101000) && ({row_reg, col_reg}<19'b1010000011001111000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010000011001111000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1010000011001111001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010000011001111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1010000011001111011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b1010000011001111100) && ({row_reg, col_reg}<19'b1010000011001111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1010000011001111110)) color_data = 12'b110111011101;

		if(({row_reg, col_reg}>=19'b1010000011001111111) && ({row_reg, col_reg}<19'b1010000100010100000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1010000100010100000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=19'b1010000100010100001) && ({row_reg, col_reg}<19'b1010000100010100011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010000100010100011) && ({row_reg, col_reg}<19'b1010000100010100101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010000100010100101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1010000100010100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010000100010100111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010000100010101000) && ({row_reg, col_reg}<19'b1010000101001111000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b1010000101001111000) && ({row_reg, col_reg}<19'b1010000101001111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010000101001111010) && ({row_reg, col_reg}<19'b1010000101001111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010000101001111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1010000101001111101)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1010000101001111110)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1010000101001111111) && ({row_reg, col_reg}<19'b1010000110010100000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1010000110010100000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=19'b1010000110010100001) && ({row_reg, col_reg}<19'b1010000110010100101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010000110010100101) && ({row_reg, col_reg}<19'b1010000110010100111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010000110010100111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010000110010101000) && ({row_reg, col_reg}<19'b1010000111001111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010000111001111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1010000111001111101)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1010000111001111110)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1010000111001111111) && ({row_reg, col_reg}<19'b1010001000010100000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1010001000010100000)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b1010001000010100001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1010001000010100010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b1010001000010100011) && ({row_reg, col_reg}<19'b1010001000010100110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1010001000010100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010001000010100111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010001000010101000) && ({row_reg, col_reg}<19'b1010001001001111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010001001001111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1010001001001111101)) color_data = 12'b101110111011;

		if(({row_reg, col_reg}>=19'b1010001001001111110) && ({row_reg, col_reg}<19'b1010001010010100000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1010001010010100000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b1010001010010100001)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1010001010010100010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010001010010100011) && ({row_reg, col_reg}<19'b1010001010010100101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b1010001010010100101) && ({row_reg, col_reg}<19'b1010001010010100111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010001010010100111) && ({row_reg, col_reg}<19'b1010001011001111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010001011001111100)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1010001011001111101)) color_data = 12'b110111011101;

		if(({row_reg, col_reg}>=19'b1010001011001111110) && ({row_reg, col_reg}<19'b1010001100010100001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1010001100010100001)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b1010001100010100010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1010001100010100011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010001100010100100) && ({row_reg, col_reg}<19'b1010001101001111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010001101001111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1010001101001111011)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1010001101001111100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=19'b1010001101001111101) && ({row_reg, col_reg}<19'b1010001110010100010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1010001110010100010)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1010001110010100011)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1010001110010100100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010001110010100101) && ({row_reg, col_reg}<19'b1010001111001111000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010001111001111000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1010001111001111001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010001111001111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1010001111001111011)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1010001111001111100)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1010001111001111101) && ({row_reg, col_reg}<19'b1010010000010100011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1010010000010100011)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1010010000010100100)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1010010000010100101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b1010010000010100110) && ({row_reg, col_reg}<19'b1010010000010110000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010010000010110000) && ({row_reg, col_reg}<19'b1010010000100111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b1010010000100111010) && ({row_reg, col_reg}<19'b1010010000100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1010010000100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b1010010000100111101) && ({row_reg, col_reg}<19'b1010010000100111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010010000100111111) && ({row_reg, col_reg}<19'b1010010000101010000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010010000101010000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1010010000101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010010000101010010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010010000101010011) && ({row_reg, col_reg}<19'b1010010000101010101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b1010010000101010101) && ({row_reg, col_reg}<19'b1010010000101010111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010010000101010111) && ({row_reg, col_reg}<19'b1010010000111001010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010010000111001010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010010000111001011) && ({row_reg, col_reg}<19'b1010010000111101001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010010000111101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010010000111101010) && ({row_reg, col_reg}<19'b1010010000111101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010010000111101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010010000111101101) && ({row_reg, col_reg}<19'b1010010000111101111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010010000111101111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010010000111110000) && ({row_reg, col_reg}<19'b1010010001001110001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b1010010001001110001) && ({row_reg, col_reg}<19'b1010010001001110011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1010010001001110011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b1010010001001110100) && ({row_reg, col_reg}<19'b1010010001001110110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010010001001110110) && ({row_reg, col_reg}<19'b1010010001001111001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010010001001111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1010010001001111010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1010010001001111011)) color_data = 12'b110111011101;

		if(({row_reg, col_reg}>=19'b1010010001001111100) && ({row_reg, col_reg}<19'b1010010010010100011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1010010010010100011)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b1010010010010100100)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1010010010010100101)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1010010010010100110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010010010010100111) && ({row_reg, col_reg}<19'b1010010010010101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010010010010101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010010010010101101) && ({row_reg, col_reg}<19'b1010010010100111000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010010010100111000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010010010100111001) && ({row_reg, col_reg}<19'b1010010010100111011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010010010100111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1010010010100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010010010100111101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010010010100111110) && ({row_reg, col_reg}<19'b1010010010101010010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b1010010010101010010) && ({row_reg, col_reg}<19'b1010010010101010101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010010010101010101) && ({row_reg, col_reg}<19'b1010010010101010111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010010010101010111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010010010101011000) && ({row_reg, col_reg}<19'b1010010010111001000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010010010111001000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010010010111001001) && ({row_reg, col_reg}<19'b1010010010111001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b1010010010111001101) && ({row_reg, col_reg}<19'b1010010010111010000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010010010111010000) && ({row_reg, col_reg}<19'b1010010010111101001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b1010010010111101001) && ({row_reg, col_reg}<19'b1010010010111101101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010010010111101101) && ({row_reg, col_reg}<19'b1010010011001110000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010010011001110000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010010011001110001) && ({row_reg, col_reg}<19'b1010010011001110011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b1010010011001110011) && ({row_reg, col_reg}<19'b1010010011001110101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010010011001110101) && ({row_reg, col_reg}<19'b1010010011001110111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b1010010011001110111) && ({row_reg, col_reg}<19'b1010010011001111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1010010011001111001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1010010011001111010)) color_data = 12'b110111011101;

		if(({row_reg, col_reg}>=19'b1010010011001111011) && ({row_reg, col_reg}<19'b1010010100010100100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1010010100010100100)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b1010010100010100101)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b1010010100010100110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=19'b1010010100010100111) && ({row_reg, col_reg}<19'b1010010100010101010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010010100010101010) && ({row_reg, col_reg}<19'b1010010100010101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b1010010100010101100) && ({row_reg, col_reg}<19'b1010010100100110000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010010100100110000) && ({row_reg, col_reg}<19'b1010010100100111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010010100100111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010010100100111011) && ({row_reg, col_reg}<19'b1010010100101010000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b1010010100101010000) && ({row_reg, col_reg}<19'b1010010100101010100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010010100101010100) && ({row_reg, col_reg}<19'b1010010100101011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b1010010100101011000) && ({row_reg, col_reg}<19'b1010010100111001001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010010100111001001) && ({row_reg, col_reg}<19'b1010010100111001011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b1010010100111001011) && ({row_reg, col_reg}<19'b1010010100111001101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010010100111001101) && ({row_reg, col_reg}<19'b1010010100111101001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b1010010100111101001) && ({row_reg, col_reg}<19'b1010010100111101011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1010010100111101011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010010100111101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1010010100111101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010010100111101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1010010100111101111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b1010010100111110000) && ({row_reg, col_reg}<19'b1010010101001110000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010010101001110000) && ({row_reg, col_reg}<19'b1010010101001110011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010010101001110011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010010101001110100) && ({row_reg, col_reg}<19'b1010010101001110110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010010101001110110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1010010101001110111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1010010101001111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1010010101001111001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1010010101001111010) && ({row_reg, col_reg}<19'b1010010110010100110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1010010110010100110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b1010010110010100111)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=19'b1010010110010101000) && ({row_reg, col_reg}<19'b1010010110010101010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=19'b1010010110010101010) && ({row_reg, col_reg}<19'b1010010110010101101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010010110010101101) && ({row_reg, col_reg}<19'b1010010110010101111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010010110010101111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010010110010110000) && ({row_reg, col_reg}<19'b1010010110100111000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010010110100111000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1010010110100111001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010010110100111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010010110100111011) && ({row_reg, col_reg}<19'b1010010110100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b1010010110100111101) && ({row_reg, col_reg}<19'b1010010110100111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010010110100111111) && ({row_reg, col_reg}<19'b1010010110101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010010110101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1010010110101010010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010010110101010011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1010010110101010100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b1010010110101010101) && ({row_reg, col_reg}<19'b1010010110101010111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010010110101010111) && ({row_reg, col_reg}<19'b1010010110111001000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010010110111001000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010010110111001001) && ({row_reg, col_reg}<19'b1010010110111001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010010110111001101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1010010110111001110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010010110111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010010110111010000) && ({row_reg, col_reg}<19'b1010010110111101001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010010110111101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010010110111101010) && ({row_reg, col_reg}<19'b1010010110111101110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010010110111101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010010110111101111) && ({row_reg, col_reg}<19'b1010010111001110000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b1010010111001110000) && ({row_reg, col_reg}<19'b1010010111001110101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1010010111001110101)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1010010111001110110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1010010111001110111)) color_data = 12'b110111011101;

		if(({row_reg, col_reg}>=19'b1010010111001111000) && ({row_reg, col_reg}<19'b1010011000010101000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1010011000010101000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b1010011000010101001)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b1010011000010101010)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1010011000010101011)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=19'b1010011000010101100) && ({row_reg, col_reg}<19'b1010011000010101110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1010011000010101110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=19'b1010011000010101111) && ({row_reg, col_reg}<19'b1010011000100111000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1010011000100111000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=19'b1010011000100111001) && ({row_reg, col_reg}<19'b1010011000100111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010011000100111011) && ({row_reg, col_reg}<19'b1010011000100111111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010011000100111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010011000101000000) && ({row_reg, col_reg}<19'b1010011000101010010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010011000101010010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1010011000101010011)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=19'b1010011000101010100) && ({row_reg, col_reg}<19'b1010011000101010111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1010011000101010111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=19'b1010011000101011000) && ({row_reg, col_reg}<19'b1010011000111001000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=19'b1010011000111001000) && ({row_reg, col_reg}<19'b1010011000111001010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1010011000111001010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=19'b1010011000111001011) && ({row_reg, col_reg}<19'b1010011000111001101)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1010011000111001101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=19'b1010011000111001110) && ({row_reg, col_reg}<19'b1010011000111010000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010011000111010000) && ({row_reg, col_reg}<19'b1010011000111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010011000111101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1010011000111101001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1010011000111101010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1010011000111101011)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1010011000111101100)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=19'b1010011000111101101) && ({row_reg, col_reg}<19'b1010011000111101111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1010011000111101111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=19'b1010011000111110000) && ({row_reg, col_reg}<19'b1010011001001110000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1010011001001110000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1010011001001110001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1010011001001110010)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1010011001001110011)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=19'b1010011001001110100) && ({row_reg, col_reg}<19'b1010011001001110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b1010011001001110110)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1010011001001110111) && ({row_reg, col_reg}<19'b1010011010010101110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=19'b1010011010010101110) && ({row_reg, col_reg}<19'b1010011010100111000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b1010011010100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1010011010100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010011010100111010) && ({row_reg, col_reg}<19'b1010011010100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010011010100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010011010100111101) && ({row_reg, col_reg}<19'b1010011010100111111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010011010100111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010011010101000000) && ({row_reg, col_reg}<19'b1010011010101010000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b1010011010101010000) && ({row_reg, col_reg}<19'b1010011010101010010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1010011010101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1010011010101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1010011010101010100) && ({row_reg, col_reg}<19'b1010011010111001110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b1010011010111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1010011010111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010011010111010000) && ({row_reg, col_reg}<19'b1010011010111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010011010111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1010011010111101001)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b1010011010111101010)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b1010011010111101011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=19'b1010011010111101100) && ({row_reg, col_reg}<19'b1010011011001110000)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1010011011001110000) && ({row_reg, col_reg}<19'b1010011100100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1010011100100111000)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b1010011100100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010011100100111010) && ({row_reg, col_reg}<19'b1010011100100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010011100100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010011100100111101) && ({row_reg, col_reg}<19'b1010011100101010010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010011100101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1010011100101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1010011100101010100) && ({row_reg, col_reg}<19'b1010011100111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1010011100111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1010011100111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010011100111010000) && ({row_reg, col_reg}<19'b1010011100111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010011100111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1010011100111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1010011100111101010) && ({row_reg, col_reg}<19'b1010011110100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1010011110100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=19'b1010011110100111001) && ({row_reg, col_reg}<19'b1010011110100111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010011110100111011) && ({row_reg, col_reg}<19'b1010011110100111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010011110100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010011110100111111) && ({row_reg, col_reg}<19'b1010011110101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010011110101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1010011110101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1010011110101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1010011110101010100) && ({row_reg, col_reg}<19'b1010011110111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1010011110111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1010011110111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010011110111010000) && ({row_reg, col_reg}<19'b1010011110111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010011110111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1010011110111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1010011110111101010) && ({row_reg, col_reg}<19'b1010100000100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1010100000100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1010100000100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010100000100111010) && ({row_reg, col_reg}<19'b1010100000100111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010100000100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010100000100111111) && ({row_reg, col_reg}<19'b1010100000101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010100000101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1010100000101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1010100000101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1010100000101010100) && ({row_reg, col_reg}<19'b1010100000111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1010100000111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1010100000111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010100000111010000) && ({row_reg, col_reg}<19'b1010100000111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010100000111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1010100000111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1010100000111101010) && ({row_reg, col_reg}<19'b1010100010100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1010100010100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1010100010100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010100010100111010) && ({row_reg, col_reg}<19'b1010100010100111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010100010100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010100010100111111) && ({row_reg, col_reg}<19'b1010100010101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010100010101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1010100010101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1010100010101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1010100010101010100) && ({row_reg, col_reg}<19'b1010100010111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1010100010111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1010100010111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010100010111010000) && ({row_reg, col_reg}<19'b1010100010111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010100010111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1010100010111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1010100010111101010) && ({row_reg, col_reg}<19'b1010100100100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1010100100100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1010100100100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010100100100111010) && ({row_reg, col_reg}<19'b1010100100100111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010100100100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010100100100111111) && ({row_reg, col_reg}<19'b1010100100101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010100100101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1010100100101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1010100100101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1010100100101010100) && ({row_reg, col_reg}<19'b1010100100111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1010100100111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1010100100111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010100100111010000) && ({row_reg, col_reg}<19'b1010100100111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010100100111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1010100100111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1010100100111101010) && ({row_reg, col_reg}<19'b1010100110100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1010100110100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1010100110100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010100110100111010) && ({row_reg, col_reg}<19'b1010100110100111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010100110100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010100110100111111) && ({row_reg, col_reg}<19'b1010100110101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010100110101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1010100110101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1010100110101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1010100110101010100) && ({row_reg, col_reg}<19'b1010100110111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1010100110111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1010100110111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010100110111010000) && ({row_reg, col_reg}<19'b1010100110111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010100110111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1010100110111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1010100110111101010) && ({row_reg, col_reg}<19'b1010101000100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1010101000100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1010101000100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010101000100111010) && ({row_reg, col_reg}<19'b1010101000100111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010101000100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010101000100111111) && ({row_reg, col_reg}<19'b1010101000101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010101000101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1010101000101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1010101000101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1010101000101010100) && ({row_reg, col_reg}<19'b1010101000111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1010101000111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1010101000111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010101000111010000) && ({row_reg, col_reg}<19'b1010101000111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010101000111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1010101000111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1010101000111101010) && ({row_reg, col_reg}<19'b1010101010100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1010101010100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1010101010100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010101010100111010) && ({row_reg, col_reg}<19'b1010101010100111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010101010100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010101010100111111) && ({row_reg, col_reg}<19'b1010101010101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010101010101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1010101010101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1010101010101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1010101010101010100) && ({row_reg, col_reg}<19'b1010101010111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1010101010111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1010101010111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010101010111010000) && ({row_reg, col_reg}<19'b1010101010111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010101010111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1010101010111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1010101010111101010) && ({row_reg, col_reg}<19'b1010101100100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1010101100100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1010101100100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010101100100111010) && ({row_reg, col_reg}<19'b1010101100100111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010101100100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010101100100111111) && ({row_reg, col_reg}<19'b1010101100101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010101100101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1010101100101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1010101100101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1010101100101010100) && ({row_reg, col_reg}<19'b1010101100111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1010101100111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1010101100111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010101100111010000) && ({row_reg, col_reg}<19'b1010101100111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010101100111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1010101100111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1010101100111101010) && ({row_reg, col_reg}<19'b1010101110100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1010101110100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1010101110100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010101110100111010) && ({row_reg, col_reg}<19'b1010101110100111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010101110100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010101110100111111) && ({row_reg, col_reg}<19'b1010101110101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010101110101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1010101110101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1010101110101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1010101110101010100) && ({row_reg, col_reg}<19'b1010101110111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1010101110111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1010101110111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010101110111010000) && ({row_reg, col_reg}<19'b1010101110111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010101110111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1010101110111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1010101110111101010) && ({row_reg, col_reg}<19'b1010110000100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1010110000100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1010110000100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010110000100111010) && ({row_reg, col_reg}<19'b1010110000100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010110000100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1010110000100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010110000100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010110000100111111) && ({row_reg, col_reg}<19'b1010110000101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010110000101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1010110000101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1010110000101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1010110000101010100) && ({row_reg, col_reg}<19'b1010110000111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1010110000111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1010110000111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010110000111010000) && ({row_reg, col_reg}<19'b1010110000111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010110000111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1010110000111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1010110000111101010) && ({row_reg, col_reg}<19'b1010110010100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1010110010100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1010110010100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010110010100111010) && ({row_reg, col_reg}<19'b1010110010100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010110010100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1010110010100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010110010100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010110010100111111) && ({row_reg, col_reg}<19'b1010110010101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010110010101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1010110010101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1010110010101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1010110010101010100) && ({row_reg, col_reg}<19'b1010110010111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1010110010111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1010110010111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010110010111010000) && ({row_reg, col_reg}<19'b1010110010111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010110010111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1010110010111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1010110010111101010) && ({row_reg, col_reg}<19'b1010110100100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1010110100100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1010110100100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010110100100111010) && ({row_reg, col_reg}<19'b1010110100100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010110100100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1010110100100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010110100100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010110100100111111) && ({row_reg, col_reg}<19'b1010110100101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010110100101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1010110100101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1010110100101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1010110100101010100) && ({row_reg, col_reg}<19'b1010110100111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1010110100111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1010110100111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010110100111010000) && ({row_reg, col_reg}<19'b1010110100111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010110100111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1010110100111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1010110100111101010) && ({row_reg, col_reg}<19'b1010110110100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1010110110100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1010110110100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010110110100111010) && ({row_reg, col_reg}<19'b1010110110100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010110110100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1010110110100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010110110100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010110110100111111) && ({row_reg, col_reg}<19'b1010110110101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010110110101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1010110110101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1010110110101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1010110110101010100) && ({row_reg, col_reg}<19'b1010110110111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1010110110111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1010110110111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010110110111010000) && ({row_reg, col_reg}<19'b1010110110111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010110110111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1010110110111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1010110110111101010) && ({row_reg, col_reg}<19'b1010111000100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1010111000100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1010111000100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010111000100111010) && ({row_reg, col_reg}<19'b1010111000100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010111000100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1010111000100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010111000100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010111000100111111) && ({row_reg, col_reg}<19'b1010111000101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010111000101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1010111000101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1010111000101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1010111000101010100) && ({row_reg, col_reg}<19'b1010111000111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1010111000111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1010111000111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010111000111010000) && ({row_reg, col_reg}<19'b1010111000111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010111000111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1010111000111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1010111000111101010) && ({row_reg, col_reg}<19'b1010111010100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1010111010100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1010111010100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010111010100111010) && ({row_reg, col_reg}<19'b1010111010100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010111010100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1010111010100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010111010100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010111010100111111) && ({row_reg, col_reg}<19'b1010111010101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010111010101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1010111010101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1010111010101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1010111010101010100) && ({row_reg, col_reg}<19'b1010111010111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1010111010111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1010111010111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010111010111010000) && ({row_reg, col_reg}<19'b1010111010111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010111010111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1010111010111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1010111010111101010) && ({row_reg, col_reg}<19'b1010111100100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1010111100100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1010111100100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010111100100111010) && ({row_reg, col_reg}<19'b1010111100100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010111100100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1010111100100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010111100100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010111100100111111) && ({row_reg, col_reg}<19'b1010111100101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010111100101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1010111100101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1010111100101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1010111100101010100) && ({row_reg, col_reg}<19'b1010111100111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1010111100111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1010111100111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010111100111010000) && ({row_reg, col_reg}<19'b1010111100111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010111100111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1010111100111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1010111100111101010) && ({row_reg, col_reg}<19'b1010111110100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1010111110100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1010111110100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010111110100111010) && ({row_reg, col_reg}<19'b1010111110100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010111110100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1010111110100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010111110100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010111110100111111) && ({row_reg, col_reg}<19'b1010111110101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010111110101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1010111110101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1010111110101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1010111110101010100) && ({row_reg, col_reg}<19'b1010111110111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1010111110111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1010111110111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1010111110111010000) && ({row_reg, col_reg}<19'b1010111110111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1010111110111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1010111110111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1010111110111101010) && ({row_reg, col_reg}<19'b1011000000100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1011000000100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1011000000100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1011000000100111010) && ({row_reg, col_reg}<19'b1011000000100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011000000100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1011000000100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011000000100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1011000000100111111) && ({row_reg, col_reg}<19'b1011000000101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011000000101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1011000000101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1011000000101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1011000000101010100) && ({row_reg, col_reg}<19'b1011000000111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1011000000111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1011000000111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1011000000111010000) && ({row_reg, col_reg}<19'b1011000000111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011000000111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1011000000111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1011000000111101010) && ({row_reg, col_reg}<19'b1011000010100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1011000010100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1011000010100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1011000010100111010) && ({row_reg, col_reg}<19'b1011000010100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011000010100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1011000010100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011000010100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1011000010100111111) && ({row_reg, col_reg}<19'b1011000010101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011000010101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1011000010101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1011000010101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1011000010101010100) && ({row_reg, col_reg}<19'b1011000010111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1011000010111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1011000010111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1011000010111010000) && ({row_reg, col_reg}<19'b1011000010111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011000010111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1011000010111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1011000010111101010) && ({row_reg, col_reg}<19'b1011000100100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1011000100100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1011000100100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1011000100100111010) && ({row_reg, col_reg}<19'b1011000100100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011000100100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1011000100100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011000100100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1011000100100111111) && ({row_reg, col_reg}<19'b1011000100101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011000100101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1011000100101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1011000100101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1011000100101010100) && ({row_reg, col_reg}<19'b1011000100111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1011000100111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1011000100111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1011000100111010000) && ({row_reg, col_reg}<19'b1011000100111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011000100111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1011000100111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1011000100111101010) && ({row_reg, col_reg}<19'b1011000110100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1011000110100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1011000110100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1011000110100111010) && ({row_reg, col_reg}<19'b1011000110100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011000110100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1011000110100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011000110100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1011000110100111111) && ({row_reg, col_reg}<19'b1011000110101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011000110101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1011000110101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1011000110101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1011000110101010100) && ({row_reg, col_reg}<19'b1011000110111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1011000110111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1011000110111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1011000110111010000) && ({row_reg, col_reg}<19'b1011000110111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011000110111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1011000110111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1011000110111101010) && ({row_reg, col_reg}<19'b1011001000100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1011001000100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1011001000100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1011001000100111010) && ({row_reg, col_reg}<19'b1011001000100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011001000100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1011001000100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011001000100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1011001000100111111) && ({row_reg, col_reg}<19'b1011001000101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011001000101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1011001000101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1011001000101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1011001000101010100) && ({row_reg, col_reg}<19'b1011001000111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1011001000111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1011001000111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1011001000111010000) && ({row_reg, col_reg}<19'b1011001000111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011001000111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1011001000111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1011001000111101010) && ({row_reg, col_reg}<19'b1011001010100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1011001010100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1011001010100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1011001010100111010) && ({row_reg, col_reg}<19'b1011001010100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011001010100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1011001010100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011001010100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1011001010100111111) && ({row_reg, col_reg}<19'b1011001010101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011001010101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1011001010101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1011001010101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1011001010101010100) && ({row_reg, col_reg}<19'b1011001010111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1011001010111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1011001010111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1011001010111010000) && ({row_reg, col_reg}<19'b1011001010111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011001010111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1011001010111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1011001010111101010) && ({row_reg, col_reg}<19'b1011001100100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1011001100100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1011001100100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1011001100100111010) && ({row_reg, col_reg}<19'b1011001100100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011001100100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1011001100100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011001100100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1011001100100111111) && ({row_reg, col_reg}<19'b1011001100101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011001100101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1011001100101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1011001100101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1011001100101010100) && ({row_reg, col_reg}<19'b1011001100111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1011001100111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1011001100111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1011001100111010000) && ({row_reg, col_reg}<19'b1011001100111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011001100111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1011001100111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1011001100111101010) && ({row_reg, col_reg}<19'b1011001110100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1011001110100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1011001110100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1011001110100111010) && ({row_reg, col_reg}<19'b1011001110100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011001110100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1011001110100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011001110100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1011001110100111111) && ({row_reg, col_reg}<19'b1011001110101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011001110101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1011001110101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1011001110101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1011001110101010100) && ({row_reg, col_reg}<19'b1011001110111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1011001110111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1011001110111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1011001110111010000) && ({row_reg, col_reg}<19'b1011001110111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011001110111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1011001110111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1011001110111101010) && ({row_reg, col_reg}<19'b1011010000100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1011010000100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1011010000100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1011010000100111010) && ({row_reg, col_reg}<19'b1011010000100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011010000100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1011010000100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011010000100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1011010000100111111) && ({row_reg, col_reg}<19'b1011010000101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011010000101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1011010000101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1011010000101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1011010000101010100) && ({row_reg, col_reg}<19'b1011010000111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1011010000111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1011010000111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1011010000111010000) && ({row_reg, col_reg}<19'b1011010000111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011010000111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1011010000111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1011010000111101010) && ({row_reg, col_reg}<19'b1011010010100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1011010010100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1011010010100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1011010010100111010) && ({row_reg, col_reg}<19'b1011010010100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011010010100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1011010010100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011010010100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1011010010100111111) && ({row_reg, col_reg}<19'b1011010010101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011010010101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1011010010101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1011010010101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1011010010101010100) && ({row_reg, col_reg}<19'b1011010010111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1011010010111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1011010010111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1011010010111010000) && ({row_reg, col_reg}<19'b1011010010111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011010010111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1011010010111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1011010010111101010) && ({row_reg, col_reg}<19'b1011010100100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1011010100100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1011010100100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1011010100100111010) && ({row_reg, col_reg}<19'b1011010100100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011010100100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1011010100100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011010100100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1011010100100111111) && ({row_reg, col_reg}<19'b1011010100101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011010100101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1011010100101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1011010100101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1011010100101010100) && ({row_reg, col_reg}<19'b1011010100111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1011010100111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1011010100111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1011010100111010000) && ({row_reg, col_reg}<19'b1011010100111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011010100111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1011010100111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1011010100111101010) && ({row_reg, col_reg}<19'b1011010110100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1011010110100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1011010110100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1011010110100111010) && ({row_reg, col_reg}<19'b1011010110100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011010110100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1011010110100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011010110100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1011010110100111111) && ({row_reg, col_reg}<19'b1011010110101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011010110101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1011010110101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1011010110101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1011010110101010100) && ({row_reg, col_reg}<19'b1011010110111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1011010110111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1011010110111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1011010110111010000) && ({row_reg, col_reg}<19'b1011010110111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011010110111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1011010110111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1011010110111101010) && ({row_reg, col_reg}<19'b1011011000100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1011011000100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1011011000100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1011011000100111010) && ({row_reg, col_reg}<19'b1011011000100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011011000100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1011011000100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011011000100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1011011000100111111) && ({row_reg, col_reg}<19'b1011011000101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011011000101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1011011000101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1011011000101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1011011000101010100) && ({row_reg, col_reg}<19'b1011011000111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1011011000111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1011011000111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1011011000111010000) && ({row_reg, col_reg}<19'b1011011000111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011011000111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1011011000111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1011011000111101010) && ({row_reg, col_reg}<19'b1011011010100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1011011010100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1011011010100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1011011010100111010) && ({row_reg, col_reg}<19'b1011011010100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011011010100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1011011010100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011011010100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1011011010100111111) && ({row_reg, col_reg}<19'b1011011010101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011011010101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1011011010101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1011011010101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1011011010101010100) && ({row_reg, col_reg}<19'b1011011010111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1011011010111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1011011010111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1011011010111010000) && ({row_reg, col_reg}<19'b1011011010111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011011010111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1011011010111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1011011010111101010) && ({row_reg, col_reg}<19'b1011011100100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1011011100100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1011011100100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1011011100100111010) && ({row_reg, col_reg}<19'b1011011100100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011011100100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1011011100100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011011100100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1011011100100111111) && ({row_reg, col_reg}<19'b1011011100101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011011100101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1011011100101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1011011100101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1011011100101010100) && ({row_reg, col_reg}<19'b1011011100111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1011011100111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1011011100111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1011011100111010000) && ({row_reg, col_reg}<19'b1011011100111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011011100111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1011011100111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1011011100111101010) && ({row_reg, col_reg}<19'b1011011110100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1011011110100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1011011110100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1011011110100111010) && ({row_reg, col_reg}<19'b1011011110100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011011110100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1011011110100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011011110100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1011011110100111111) && ({row_reg, col_reg}<19'b1011011110101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011011110101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1011011110101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1011011110101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1011011110101010100) && ({row_reg, col_reg}<19'b1011011110111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1011011110111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1011011110111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1011011110111010000) && ({row_reg, col_reg}<19'b1011011110111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011011110111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1011011110111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1011011110111101010) && ({row_reg, col_reg}<19'b1011100000100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1011100000100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1011100000100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1011100000100111010) && ({row_reg, col_reg}<19'b1011100000100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011100000100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1011100000100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011100000100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1011100000100111111) && ({row_reg, col_reg}<19'b1011100000101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011100000101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1011100000101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1011100000101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1011100000101010100) && ({row_reg, col_reg}<19'b1011100000111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1011100000111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1011100000111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1011100000111010000) && ({row_reg, col_reg}<19'b1011100000111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011100000111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1011100000111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1011100000111101010) && ({row_reg, col_reg}<19'b1011100010100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1011100010100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1011100010100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1011100010100111010) && ({row_reg, col_reg}<19'b1011100010100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011100010100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1011100010100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011100010100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1011100010100111111) && ({row_reg, col_reg}<19'b1011100010101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011100010101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1011100010101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1011100010101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1011100010101010100) && ({row_reg, col_reg}<19'b1011100010111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1011100010111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1011100010111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1011100010111010000) && ({row_reg, col_reg}<19'b1011100010111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011100010111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1011100010111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1011100010111101010) && ({row_reg, col_reg}<19'b1011100100100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1011100100100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1011100100100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1011100100100111010) && ({row_reg, col_reg}<19'b1011100100100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011100100100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1011100100100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011100100100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1011100100100111111) && ({row_reg, col_reg}<19'b1011100100101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011100100101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1011100100101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1011100100101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1011100100101010100) && ({row_reg, col_reg}<19'b1011100100111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1011100100111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1011100100111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1011100100111010000) && ({row_reg, col_reg}<19'b1011100100111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011100100111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1011100100111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1011100100111101010) && ({row_reg, col_reg}<19'b1011100110100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1011100110100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1011100110100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1011100110100111010) && ({row_reg, col_reg}<19'b1011100110100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011100110100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1011100110100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011100110100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1011100110100111111) && ({row_reg, col_reg}<19'b1011100110101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011100110101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1011100110101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1011100110101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1011100110101010100) && ({row_reg, col_reg}<19'b1011100110111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1011100110111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1011100110111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1011100110111010000) && ({row_reg, col_reg}<19'b1011100110111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011100110111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1011100110111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1011100110111101010) && ({row_reg, col_reg}<19'b1011101000100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1011101000100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1011101000100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1011101000100111010) && ({row_reg, col_reg}<19'b1011101000100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011101000100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1011101000100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011101000100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1011101000100111111) && ({row_reg, col_reg}<19'b1011101000101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011101000101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1011101000101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1011101000101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1011101000101010100) && ({row_reg, col_reg}<19'b1011101000111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1011101000111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1011101000111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1011101000111010000) && ({row_reg, col_reg}<19'b1011101000111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011101000111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1011101000111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1011101000111101010) && ({row_reg, col_reg}<19'b1011101010100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1011101010100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1011101010100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1011101010100111010) && ({row_reg, col_reg}<19'b1011101010100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011101010100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1011101010100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011101010100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1011101010100111111) && ({row_reg, col_reg}<19'b1011101010101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011101010101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1011101010101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1011101010101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1011101010101010100) && ({row_reg, col_reg}<19'b1011101010111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1011101010111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1011101010111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1011101010111010000) && ({row_reg, col_reg}<19'b1011101010111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011101010111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1011101010111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1011101010111101010) && ({row_reg, col_reg}<19'b1011101100100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1011101100100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1011101100100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1011101100100111010) && ({row_reg, col_reg}<19'b1011101100100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011101100100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1011101100100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011101100100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1011101100100111111) && ({row_reg, col_reg}<19'b1011101100101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011101100101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1011101100101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1011101100101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1011101100101010100) && ({row_reg, col_reg}<19'b1011101100111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1011101100111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1011101100111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1011101100111010000) && ({row_reg, col_reg}<19'b1011101100111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011101100111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1011101100111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1011101100111101010) && ({row_reg, col_reg}<19'b1011101110100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1011101110100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1011101110100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1011101110100111010) && ({row_reg, col_reg}<19'b1011101110100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011101110100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1011101110100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011101110100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1011101110100111111) && ({row_reg, col_reg}<19'b1011101110101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011101110101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1011101110101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1011101110101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1011101110101010100) && ({row_reg, col_reg}<19'b1011101110111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1011101110111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1011101110111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1011101110111010000) && ({row_reg, col_reg}<19'b1011101110111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011101110111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1011101110111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1011101110111101010) && ({row_reg, col_reg}<19'b1011110000100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1011110000100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1011110000100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1011110000100111010) && ({row_reg, col_reg}<19'b1011110000100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011110000100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1011110000100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011110000100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1011110000100111111) && ({row_reg, col_reg}<19'b1011110000101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011110000101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1011110000101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1011110000101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1011110000101010100) && ({row_reg, col_reg}<19'b1011110000111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1011110000111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1011110000111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1011110000111010000) && ({row_reg, col_reg}<19'b1011110000111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011110000111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1011110000111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1011110000111101010) && ({row_reg, col_reg}<19'b1011110010100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1011110010100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1011110010100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1011110010100111010) && ({row_reg, col_reg}<19'b1011110010100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011110010100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1011110010100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011110010100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1011110010100111111) && ({row_reg, col_reg}<19'b1011110010101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011110010101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1011110010101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1011110010101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1011110010101010100) && ({row_reg, col_reg}<19'b1011110010111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1011110010111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1011110010111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1011110010111010000) && ({row_reg, col_reg}<19'b1011110010111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011110010111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1011110010111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1011110010111101010) && ({row_reg, col_reg}<19'b1011110100100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1011110100100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1011110100100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1011110100100111010) && ({row_reg, col_reg}<19'b1011110100100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011110100100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1011110100100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011110100100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1011110100100111111) && ({row_reg, col_reg}<19'b1011110100101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011110100101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1011110100101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1011110100101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1011110100101010100) && ({row_reg, col_reg}<19'b1011110100111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1011110100111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1011110100111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1011110100111010000) && ({row_reg, col_reg}<19'b1011110100111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011110100111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1011110100111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1011110100111101010) && ({row_reg, col_reg}<19'b1011110110100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1011110110100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1011110110100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1011110110100111010) && ({row_reg, col_reg}<19'b1011110110100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011110110100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1011110110100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011110110100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1011110110100111111) && ({row_reg, col_reg}<19'b1011110110101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011110110101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1011110110101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1011110110101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1011110110101010100) && ({row_reg, col_reg}<19'b1011110110111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1011110110111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1011110110111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1011110110111010000) && ({row_reg, col_reg}<19'b1011110110111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011110110111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1011110110111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1011110110111101010) && ({row_reg, col_reg}<19'b1011111000100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1011111000100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1011111000100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1011111000100111010) && ({row_reg, col_reg}<19'b1011111000100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011111000100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1011111000100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011111000100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1011111000100111111) && ({row_reg, col_reg}<19'b1011111000101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011111000101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1011111000101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1011111000101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1011111000101010100) && ({row_reg, col_reg}<19'b1011111000111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1011111000111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1011111000111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1011111000111010000) && ({row_reg, col_reg}<19'b1011111000111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011111000111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1011111000111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1011111000111101010) && ({row_reg, col_reg}<19'b1011111010100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1011111010100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1011111010100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1011111010100111010) && ({row_reg, col_reg}<19'b1011111010100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011111010100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1011111010100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011111010100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1011111010100111111) && ({row_reg, col_reg}<19'b1011111010101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011111010101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1011111010101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1011111010101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1011111010101010100) && ({row_reg, col_reg}<19'b1011111010111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1011111010111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1011111010111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1011111010111010000) && ({row_reg, col_reg}<19'b1011111010111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011111010111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1011111010111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1011111010111101010) && ({row_reg, col_reg}<19'b1011111100100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1011111100100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1011111100100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1011111100100111010) && ({row_reg, col_reg}<19'b1011111100100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011111100100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1011111100100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011111100100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1011111100100111111) && ({row_reg, col_reg}<19'b1011111100101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011111100101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1011111100101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1011111100101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1011111100101010100) && ({row_reg, col_reg}<19'b1011111100111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1011111100111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1011111100111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1011111100111010000) && ({row_reg, col_reg}<19'b1011111100111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011111100111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1011111100111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1011111100111101010) && ({row_reg, col_reg}<19'b1011111110100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1011111110100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1011111110100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1011111110100111010) && ({row_reg, col_reg}<19'b1011111110100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011111110100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1011111110100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011111110100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1011111110100111111) && ({row_reg, col_reg}<19'b1011111110101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011111110101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1011111110101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1011111110101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1011111110101010100) && ({row_reg, col_reg}<19'b1011111110111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1011111110111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1011111110111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1011111110111010000) && ({row_reg, col_reg}<19'b1011111110111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1011111110111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1011111110111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1011111110111101010) && ({row_reg, col_reg}<19'b1100000000100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1100000000100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1100000000100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1100000000100111010) && ({row_reg, col_reg}<19'b1100000000100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100000000100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1100000000100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100000000100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1100000000100111111) && ({row_reg, col_reg}<19'b1100000000101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100000000101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1100000000101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1100000000101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1100000000101010100) && ({row_reg, col_reg}<19'b1100000000111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1100000000111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1100000000111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1100000000111010000) && ({row_reg, col_reg}<19'b1100000000111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100000000111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1100000000111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1100000000111101010) && ({row_reg, col_reg}<19'b1100000010100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1100000010100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1100000010100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1100000010100111010) && ({row_reg, col_reg}<19'b1100000010100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100000010100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1100000010100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100000010100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1100000010100111111) && ({row_reg, col_reg}<19'b1100000010101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100000010101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1100000010101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1100000010101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1100000010101010100) && ({row_reg, col_reg}<19'b1100000010111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1100000010111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1100000010111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1100000010111010000) && ({row_reg, col_reg}<19'b1100000010111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100000010111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1100000010111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1100000010111101010) && ({row_reg, col_reg}<19'b1100000100100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1100000100100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1100000100100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1100000100100111010) && ({row_reg, col_reg}<19'b1100000100100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100000100100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1100000100100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100000100100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1100000100100111111) && ({row_reg, col_reg}<19'b1100000100101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100000100101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1100000100101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1100000100101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1100000100101010100) && ({row_reg, col_reg}<19'b1100000100111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1100000100111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1100000100111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1100000100111010000) && ({row_reg, col_reg}<19'b1100000100111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100000100111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1100000100111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1100000100111101010) && ({row_reg, col_reg}<19'b1100000110100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1100000110100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1100000110100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1100000110100111010) && ({row_reg, col_reg}<19'b1100000110100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100000110100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1100000110100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100000110100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1100000110100111111) && ({row_reg, col_reg}<19'b1100000110101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100000110101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1100000110101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1100000110101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1100000110101010100) && ({row_reg, col_reg}<19'b1100000110111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1100000110111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1100000110111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1100000110111010000) && ({row_reg, col_reg}<19'b1100000110111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100000110111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1100000110111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1100000110111101010) && ({row_reg, col_reg}<19'b1100001000100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1100001000100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1100001000100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1100001000100111010) && ({row_reg, col_reg}<19'b1100001000100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100001000100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1100001000100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100001000100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1100001000100111111) && ({row_reg, col_reg}<19'b1100001000101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100001000101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1100001000101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1100001000101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1100001000101010100) && ({row_reg, col_reg}<19'b1100001000111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1100001000111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1100001000111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1100001000111010000) && ({row_reg, col_reg}<19'b1100001000111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100001000111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1100001000111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1100001000111101010) && ({row_reg, col_reg}<19'b1100001010100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1100001010100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1100001010100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1100001010100111010) && ({row_reg, col_reg}<19'b1100001010100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100001010100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1100001010100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100001010100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1100001010100111111) && ({row_reg, col_reg}<19'b1100001010101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100001010101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1100001010101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1100001010101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1100001010101010100) && ({row_reg, col_reg}<19'b1100001010111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1100001010111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1100001010111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1100001010111010000) && ({row_reg, col_reg}<19'b1100001010111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100001010111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1100001010111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1100001010111101010) && ({row_reg, col_reg}<19'b1100001100100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1100001100100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1100001100100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1100001100100111010) && ({row_reg, col_reg}<19'b1100001100100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100001100100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1100001100100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100001100100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1100001100100111111) && ({row_reg, col_reg}<19'b1100001100101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100001100101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1100001100101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1100001100101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1100001100101010100) && ({row_reg, col_reg}<19'b1100001100111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1100001100111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1100001100111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1100001100111010000) && ({row_reg, col_reg}<19'b1100001100111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100001100111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1100001100111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1100001100111101010) && ({row_reg, col_reg}<19'b1100001110100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1100001110100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1100001110100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1100001110100111010) && ({row_reg, col_reg}<19'b1100001110100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100001110100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1100001110100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100001110100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1100001110100111111) && ({row_reg, col_reg}<19'b1100001110101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100001110101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1100001110101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1100001110101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1100001110101010100) && ({row_reg, col_reg}<19'b1100001110111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1100001110111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1100001110111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1100001110111010000) && ({row_reg, col_reg}<19'b1100001110111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100001110111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1100001110111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1100001110111101010) && ({row_reg, col_reg}<19'b1100010000100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1100010000100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1100010000100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1100010000100111010) && ({row_reg, col_reg}<19'b1100010000100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100010000100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1100010000100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100010000100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1100010000100111111) && ({row_reg, col_reg}<19'b1100010000101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100010000101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1100010000101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1100010000101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1100010000101010100) && ({row_reg, col_reg}<19'b1100010000111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1100010000111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1100010000111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1100010000111010000) && ({row_reg, col_reg}<19'b1100010000111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100010000111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1100010000111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1100010000111101010) && ({row_reg, col_reg}<19'b1100010010100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1100010010100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1100010010100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1100010010100111010) && ({row_reg, col_reg}<19'b1100010010100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100010010100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1100010010100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100010010100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1100010010100111111) && ({row_reg, col_reg}<19'b1100010010101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100010010101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1100010010101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1100010010101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1100010010101010100) && ({row_reg, col_reg}<19'b1100010010111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1100010010111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1100010010111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1100010010111010000) && ({row_reg, col_reg}<19'b1100010010111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100010010111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1100010010111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1100010010111101010) && ({row_reg, col_reg}<19'b1100010100100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1100010100100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1100010100100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1100010100100111010) && ({row_reg, col_reg}<19'b1100010100100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100010100100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1100010100100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100010100100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1100010100100111111) && ({row_reg, col_reg}<19'b1100010100101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100010100101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1100010100101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1100010100101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1100010100101010100) && ({row_reg, col_reg}<19'b1100010100111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1100010100111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1100010100111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1100010100111010000) && ({row_reg, col_reg}<19'b1100010100111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100010100111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1100010100111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1100010100111101010) && ({row_reg, col_reg}<19'b1100010110100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1100010110100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1100010110100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1100010110100111010) && ({row_reg, col_reg}<19'b1100010110100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100010110100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1100010110100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100010110100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1100010110100111111) && ({row_reg, col_reg}<19'b1100010110101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100010110101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1100010110101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1100010110101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1100010110101010100) && ({row_reg, col_reg}<19'b1100010110111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1100010110111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1100010110111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1100010110111010000) && ({row_reg, col_reg}<19'b1100010110111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100010110111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1100010110111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1100010110111101010) && ({row_reg, col_reg}<19'b1100011000100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1100011000100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1100011000100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1100011000100111010) && ({row_reg, col_reg}<19'b1100011000100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100011000100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1100011000100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100011000100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1100011000100111111) && ({row_reg, col_reg}<19'b1100011000101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100011000101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1100011000101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1100011000101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1100011000101010100) && ({row_reg, col_reg}<19'b1100011000111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1100011000111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1100011000111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1100011000111010000) && ({row_reg, col_reg}<19'b1100011000111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100011000111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1100011000111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1100011000111101010) && ({row_reg, col_reg}<19'b1100011010100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1100011010100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1100011010100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1100011010100111010) && ({row_reg, col_reg}<19'b1100011010100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100011010100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1100011010100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100011010100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1100011010100111111) && ({row_reg, col_reg}<19'b1100011010101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100011010101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1100011010101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1100011010101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1100011010101010100) && ({row_reg, col_reg}<19'b1100011010111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1100011010111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1100011010111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1100011010111010000) && ({row_reg, col_reg}<19'b1100011010111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100011010111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1100011010111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1100011010111101010) && ({row_reg, col_reg}<19'b1100011100100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1100011100100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1100011100100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1100011100100111010) && ({row_reg, col_reg}<19'b1100011100100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100011100100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1100011100100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100011100100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1100011100100111111) && ({row_reg, col_reg}<19'b1100011100101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100011100101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1100011100101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1100011100101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1100011100101010100) && ({row_reg, col_reg}<19'b1100011100111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1100011100111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1100011100111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1100011100111010000) && ({row_reg, col_reg}<19'b1100011100111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100011100111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1100011100111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1100011100111101010) && ({row_reg, col_reg}<19'b1100011110100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1100011110100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1100011110100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1100011110100111010) && ({row_reg, col_reg}<19'b1100011110100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100011110100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1100011110100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100011110100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1100011110100111111) && ({row_reg, col_reg}<19'b1100011110101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100011110101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1100011110101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1100011110101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1100011110101010100) && ({row_reg, col_reg}<19'b1100011110111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1100011110111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1100011110111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1100011110111010000) && ({row_reg, col_reg}<19'b1100011110111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100011110111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1100011110111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1100011110111101010) && ({row_reg, col_reg}<19'b1100100000100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1100100000100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1100100000100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1100100000100111010) && ({row_reg, col_reg}<19'b1100100000100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100100000100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1100100000100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100100000100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1100100000100111111) && ({row_reg, col_reg}<19'b1100100000101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100100000101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1100100000101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1100100000101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1100100000101010100) && ({row_reg, col_reg}<19'b1100100000111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1100100000111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1100100000111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1100100000111010000) && ({row_reg, col_reg}<19'b1100100000111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100100000111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1100100000111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1100100000111101010) && ({row_reg, col_reg}<19'b1100100010100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1100100010100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1100100010100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1100100010100111010) && ({row_reg, col_reg}<19'b1100100010100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100100010100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1100100010100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100100010100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1100100010100111111) && ({row_reg, col_reg}<19'b1100100010101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100100010101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1100100010101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1100100010101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1100100010101010100) && ({row_reg, col_reg}<19'b1100100010111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1100100010111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1100100010111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1100100010111010000) && ({row_reg, col_reg}<19'b1100100010111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100100010111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1100100010111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1100100010111101010) && ({row_reg, col_reg}<19'b1100100100100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1100100100100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1100100100100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1100100100100111010) && ({row_reg, col_reg}<19'b1100100100100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100100100100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1100100100100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100100100100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1100100100100111111) && ({row_reg, col_reg}<19'b1100100100101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100100100101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1100100100101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1100100100101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1100100100101010100) && ({row_reg, col_reg}<19'b1100100100111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1100100100111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1100100100111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1100100100111010000) && ({row_reg, col_reg}<19'b1100100100111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100100100111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1100100100111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1100100100111101010) && ({row_reg, col_reg}<19'b1100100110100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1100100110100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1100100110100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1100100110100111010) && ({row_reg, col_reg}<19'b1100100110100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100100110100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1100100110100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100100110100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1100100110100111111) && ({row_reg, col_reg}<19'b1100100110101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100100110101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1100100110101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1100100110101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1100100110101010100) && ({row_reg, col_reg}<19'b1100100110111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1100100110111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1100100110111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1100100110111010000) && ({row_reg, col_reg}<19'b1100100110111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100100110111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1100100110111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1100100110111101010) && ({row_reg, col_reg}<19'b1100101000100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1100101000100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1100101000100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1100101000100111010) && ({row_reg, col_reg}<19'b1100101000100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100101000100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1100101000100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100101000100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1100101000100111111) && ({row_reg, col_reg}<19'b1100101000101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100101000101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1100101000101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1100101000101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1100101000101010100) && ({row_reg, col_reg}<19'b1100101000111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1100101000111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1100101000111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1100101000111010000) && ({row_reg, col_reg}<19'b1100101000111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100101000111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1100101000111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1100101000111101010) && ({row_reg, col_reg}<19'b1100101010100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1100101010100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1100101010100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1100101010100111010) && ({row_reg, col_reg}<19'b1100101010100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100101010100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1100101010100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100101010100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1100101010100111111) && ({row_reg, col_reg}<19'b1100101010101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100101010101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1100101010101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1100101010101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1100101010101010100) && ({row_reg, col_reg}<19'b1100101010111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1100101010111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1100101010111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1100101010111010000) && ({row_reg, col_reg}<19'b1100101010111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100101010111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1100101010111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1100101010111101010) && ({row_reg, col_reg}<19'b1100101100100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1100101100100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1100101100100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1100101100100111010) && ({row_reg, col_reg}<19'b1100101100100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100101100100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1100101100100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100101100100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1100101100100111111) && ({row_reg, col_reg}<19'b1100101100101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100101100101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1100101100101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1100101100101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1100101100101010100) && ({row_reg, col_reg}<19'b1100101100111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1100101100111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1100101100111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1100101100111010000) && ({row_reg, col_reg}<19'b1100101100111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100101100111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1100101100111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1100101100111101010) && ({row_reg, col_reg}<19'b1100101110100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1100101110100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1100101110100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1100101110100111010) && ({row_reg, col_reg}<19'b1100101110100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100101110100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1100101110100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100101110100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1100101110100111111) && ({row_reg, col_reg}<19'b1100101110101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100101110101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1100101110101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1100101110101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1100101110101010100) && ({row_reg, col_reg}<19'b1100101110111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1100101110111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1100101110111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1100101110111010000) && ({row_reg, col_reg}<19'b1100101110111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100101110111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1100101110111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1100101110111101010) && ({row_reg, col_reg}<19'b1100110000100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1100110000100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1100110000100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1100110000100111010) && ({row_reg, col_reg}<19'b1100110000100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100110000100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1100110000100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100110000100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1100110000100111111) && ({row_reg, col_reg}<19'b1100110000101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100110000101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1100110000101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1100110000101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1100110000101010100) && ({row_reg, col_reg}<19'b1100110000111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1100110000111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1100110000111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1100110000111010000) && ({row_reg, col_reg}<19'b1100110000111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100110000111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1100110000111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1100110000111101010) && ({row_reg, col_reg}<19'b1100110010100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1100110010100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1100110010100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1100110010100111010) && ({row_reg, col_reg}<19'b1100110010100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100110010100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1100110010100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100110010100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1100110010100111111) && ({row_reg, col_reg}<19'b1100110010101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100110010101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1100110010101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1100110010101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1100110010101010100) && ({row_reg, col_reg}<19'b1100110010111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1100110010111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1100110010111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1100110010111010000) && ({row_reg, col_reg}<19'b1100110010111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100110010111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1100110010111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1100110010111101010) && ({row_reg, col_reg}<19'b1100110100100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1100110100100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1100110100100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1100110100100111010) && ({row_reg, col_reg}<19'b1100110100100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100110100100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1100110100100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100110100100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1100110100100111111) && ({row_reg, col_reg}<19'b1100110100101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100110100101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1100110100101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1100110100101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1100110100101010100) && ({row_reg, col_reg}<19'b1100110100111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1100110100111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1100110100111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1100110100111010000) && ({row_reg, col_reg}<19'b1100110100111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100110100111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1100110100111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1100110100111101010) && ({row_reg, col_reg}<19'b1100110110100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1100110110100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1100110110100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1100110110100111010) && ({row_reg, col_reg}<19'b1100110110100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100110110100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1100110110100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100110110100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1100110110100111111) && ({row_reg, col_reg}<19'b1100110110101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100110110101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1100110110101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1100110110101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1100110110101010100) && ({row_reg, col_reg}<19'b1100110110111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1100110110111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1100110110111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1100110110111010000) && ({row_reg, col_reg}<19'b1100110110111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100110110111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1100110110111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1100110110111101010) && ({row_reg, col_reg}<19'b1100111000100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1100111000100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1100111000100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1100111000100111010) && ({row_reg, col_reg}<19'b1100111000100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100111000100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1100111000100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100111000100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1100111000100111111) && ({row_reg, col_reg}<19'b1100111000101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100111000101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1100111000101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1100111000101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1100111000101010100) && ({row_reg, col_reg}<19'b1100111000111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1100111000111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1100111000111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1100111000111010000) && ({row_reg, col_reg}<19'b1100111000111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100111000111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1100111000111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1100111000111101010) && ({row_reg, col_reg}<19'b1100111010100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1100111010100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1100111010100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1100111010100111010) && ({row_reg, col_reg}<19'b1100111010100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100111010100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1100111010100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100111010100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1100111010100111111) && ({row_reg, col_reg}<19'b1100111010101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100111010101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1100111010101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1100111010101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1100111010101010100) && ({row_reg, col_reg}<19'b1100111010111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1100111010111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1100111010111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1100111010111010000) && ({row_reg, col_reg}<19'b1100111010111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100111010111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1100111010111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1100111010111101010) && ({row_reg, col_reg}<19'b1100111100100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1100111100100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1100111100100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1100111100100111010) && ({row_reg, col_reg}<19'b1100111100100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100111100100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1100111100100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100111100100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1100111100100111111) && ({row_reg, col_reg}<19'b1100111100101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100111100101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1100111100101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1100111100101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1100111100101010100) && ({row_reg, col_reg}<19'b1100111100111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1100111100111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1100111100111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1100111100111010000) && ({row_reg, col_reg}<19'b1100111100111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100111100111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1100111100111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1100111100111101010) && ({row_reg, col_reg}<19'b1100111110100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1100111110100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1100111110100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1100111110100111010) && ({row_reg, col_reg}<19'b1100111110100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100111110100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1100111110100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100111110100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1100111110100111111) && ({row_reg, col_reg}<19'b1100111110101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100111110101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1100111110101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1100111110101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1100111110101010100) && ({row_reg, col_reg}<19'b1100111110111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1100111110111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1100111110111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1100111110111010000) && ({row_reg, col_reg}<19'b1100111110111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1100111110111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1100111110111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1100111110111101010) && ({row_reg, col_reg}<19'b1101000000100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1101000000100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1101000000100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1101000000100111010) && ({row_reg, col_reg}<19'b1101000000100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101000000100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1101000000100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101000000100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1101000000100111111) && ({row_reg, col_reg}<19'b1101000000101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101000000101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1101000000101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1101000000101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1101000000101010100) && ({row_reg, col_reg}<19'b1101000000111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1101000000111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1101000000111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1101000000111010000) && ({row_reg, col_reg}<19'b1101000000111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101000000111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1101000000111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1101000000111101010) && ({row_reg, col_reg}<19'b1101000010100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1101000010100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1101000010100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1101000010100111010) && ({row_reg, col_reg}<19'b1101000010100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101000010100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1101000010100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101000010100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1101000010100111111) && ({row_reg, col_reg}<19'b1101000010101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101000010101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1101000010101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1101000010101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1101000010101010100) && ({row_reg, col_reg}<19'b1101000010111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1101000010111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1101000010111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1101000010111010000) && ({row_reg, col_reg}<19'b1101000010111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101000010111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1101000010111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1101000010111101010) && ({row_reg, col_reg}<19'b1101000100100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1101000100100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1101000100100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1101000100100111010) && ({row_reg, col_reg}<19'b1101000100100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101000100100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1101000100100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101000100100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1101000100100111111) && ({row_reg, col_reg}<19'b1101000100101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101000100101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1101000100101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1101000100101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1101000100101010100) && ({row_reg, col_reg}<19'b1101000100111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1101000100111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1101000100111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1101000100111010000) && ({row_reg, col_reg}<19'b1101000100111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101000100111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1101000100111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1101000100111101010) && ({row_reg, col_reg}<19'b1101000110100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1101000110100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1101000110100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1101000110100111010) && ({row_reg, col_reg}<19'b1101000110100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101000110100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1101000110100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101000110100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1101000110100111111) && ({row_reg, col_reg}<19'b1101000110101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101000110101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1101000110101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1101000110101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1101000110101010100) && ({row_reg, col_reg}<19'b1101000110111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1101000110111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1101000110111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1101000110111010000) && ({row_reg, col_reg}<19'b1101000110111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101000110111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1101000110111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1101000110111101010) && ({row_reg, col_reg}<19'b1101001000100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1101001000100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1101001000100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1101001000100111010) && ({row_reg, col_reg}<19'b1101001000100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101001000100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1101001000100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101001000100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1101001000100111111) && ({row_reg, col_reg}<19'b1101001000101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101001000101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1101001000101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1101001000101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1101001000101010100) && ({row_reg, col_reg}<19'b1101001000111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1101001000111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1101001000111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1101001000111010000) && ({row_reg, col_reg}<19'b1101001000111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101001000111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1101001000111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1101001000111101010) && ({row_reg, col_reg}<19'b1101001010100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1101001010100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1101001010100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1101001010100111010) && ({row_reg, col_reg}<19'b1101001010100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101001010100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1101001010100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101001010100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1101001010100111111) && ({row_reg, col_reg}<19'b1101001010101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101001010101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1101001010101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1101001010101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1101001010101010100) && ({row_reg, col_reg}<19'b1101001010111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1101001010111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1101001010111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1101001010111010000) && ({row_reg, col_reg}<19'b1101001010111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101001010111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1101001010111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1101001010111101010) && ({row_reg, col_reg}<19'b1101001100100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1101001100100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1101001100100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1101001100100111010) && ({row_reg, col_reg}<19'b1101001100100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101001100100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1101001100100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101001100100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1101001100100111111) && ({row_reg, col_reg}<19'b1101001100101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101001100101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1101001100101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1101001100101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1101001100101010100) && ({row_reg, col_reg}<19'b1101001100111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1101001100111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1101001100111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1101001100111010000) && ({row_reg, col_reg}<19'b1101001100111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101001100111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1101001100111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1101001100111101010) && ({row_reg, col_reg}<19'b1101001110100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1101001110100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1101001110100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1101001110100111010) && ({row_reg, col_reg}<19'b1101001110100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101001110100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1101001110100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101001110100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1101001110100111111) && ({row_reg, col_reg}<19'b1101001110101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101001110101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1101001110101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1101001110101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1101001110101010100) && ({row_reg, col_reg}<19'b1101001110111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1101001110111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1101001110111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1101001110111010000) && ({row_reg, col_reg}<19'b1101001110111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101001110111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1101001110111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1101001110111101010) && ({row_reg, col_reg}<19'b1101010000100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1101010000100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1101010000100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1101010000100111010) && ({row_reg, col_reg}<19'b1101010000100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101010000100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1101010000100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101010000100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1101010000100111111) && ({row_reg, col_reg}<19'b1101010000101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101010000101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1101010000101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1101010000101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1101010000101010100) && ({row_reg, col_reg}<19'b1101010000111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1101010000111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1101010000111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1101010000111010000) && ({row_reg, col_reg}<19'b1101010000111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101010000111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1101010000111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1101010000111101010) && ({row_reg, col_reg}<19'b1101010010100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1101010010100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1101010010100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1101010010100111010) && ({row_reg, col_reg}<19'b1101010010100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101010010100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1101010010100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101010010100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1101010010100111111) && ({row_reg, col_reg}<19'b1101010010101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101010010101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1101010010101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1101010010101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1101010010101010100) && ({row_reg, col_reg}<19'b1101010010111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1101010010111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1101010010111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1101010010111010000) && ({row_reg, col_reg}<19'b1101010010111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101010010111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1101010010111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1101010010111101010) && ({row_reg, col_reg}<19'b1101010100100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1101010100100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1101010100100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1101010100100111010) && ({row_reg, col_reg}<19'b1101010100100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101010100100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1101010100100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101010100100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1101010100100111111) && ({row_reg, col_reg}<19'b1101010100101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101010100101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1101010100101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1101010100101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1101010100101010100) && ({row_reg, col_reg}<19'b1101010100111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1101010100111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1101010100111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1101010100111010000) && ({row_reg, col_reg}<19'b1101010100111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101010100111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1101010100111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1101010100111101010) && ({row_reg, col_reg}<19'b1101010110100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1101010110100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1101010110100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1101010110100111010) && ({row_reg, col_reg}<19'b1101010110100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101010110100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1101010110100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101010110100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1101010110100111111) && ({row_reg, col_reg}<19'b1101010110101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101010110101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1101010110101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1101010110101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1101010110101010100) && ({row_reg, col_reg}<19'b1101010110111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1101010110111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1101010110111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1101010110111010000) && ({row_reg, col_reg}<19'b1101010110111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101010110111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1101010110111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1101010110111101010) && ({row_reg, col_reg}<19'b1101011000100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1101011000100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1101011000100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1101011000100111010) && ({row_reg, col_reg}<19'b1101011000100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101011000100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1101011000100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101011000100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1101011000100111111) && ({row_reg, col_reg}<19'b1101011000101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101011000101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1101011000101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1101011000101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1101011000101010100) && ({row_reg, col_reg}<19'b1101011000111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1101011000111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1101011000111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1101011000111010000) && ({row_reg, col_reg}<19'b1101011000111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101011000111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1101011000111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1101011000111101010) && ({row_reg, col_reg}<19'b1101011010100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1101011010100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1101011010100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1101011010100111010) && ({row_reg, col_reg}<19'b1101011010100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101011010100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1101011010100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101011010100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1101011010100111111) && ({row_reg, col_reg}<19'b1101011010101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101011010101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1101011010101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1101011010101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1101011010101010100) && ({row_reg, col_reg}<19'b1101011010111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1101011010111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1101011010111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1101011010111010000) && ({row_reg, col_reg}<19'b1101011010111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101011010111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1101011010111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1101011010111101010) && ({row_reg, col_reg}<19'b1101011100100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1101011100100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1101011100100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1101011100100111010) && ({row_reg, col_reg}<19'b1101011100100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101011100100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1101011100100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101011100100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1101011100100111111) && ({row_reg, col_reg}<19'b1101011100101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101011100101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1101011100101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1101011100101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1101011100101010100) && ({row_reg, col_reg}<19'b1101011100111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1101011100111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1101011100111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1101011100111010000) && ({row_reg, col_reg}<19'b1101011100111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101011100111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1101011100111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1101011100111101010) && ({row_reg, col_reg}<19'b1101011110100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1101011110100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1101011110100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1101011110100111010) && ({row_reg, col_reg}<19'b1101011110100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101011110100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1101011110100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101011110100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1101011110100111111) && ({row_reg, col_reg}<19'b1101011110101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101011110101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1101011110101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1101011110101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1101011110101010100) && ({row_reg, col_reg}<19'b1101011110111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1101011110111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1101011110111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1101011110111010000) && ({row_reg, col_reg}<19'b1101011110111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101011110111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1101011110111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1101011110111101010) && ({row_reg, col_reg}<19'b1101100000100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1101100000100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1101100000100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1101100000100111010) && ({row_reg, col_reg}<19'b1101100000100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101100000100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1101100000100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101100000100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1101100000100111111) && ({row_reg, col_reg}<19'b1101100000101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101100000101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1101100000101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1101100000101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1101100000101010100) && ({row_reg, col_reg}<19'b1101100000111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1101100000111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1101100000111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1101100000111010000) && ({row_reg, col_reg}<19'b1101100000111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101100000111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1101100000111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1101100000111101010) && ({row_reg, col_reg}<19'b1101100010100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1101100010100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1101100010100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1101100010100111010) && ({row_reg, col_reg}<19'b1101100010100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101100010100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1101100010100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101100010100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1101100010100111111) && ({row_reg, col_reg}<19'b1101100010101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101100010101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1101100010101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1101100010101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1101100010101010100) && ({row_reg, col_reg}<19'b1101100010111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1101100010111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1101100010111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1101100010111010000) && ({row_reg, col_reg}<19'b1101100010111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101100010111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1101100010111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1101100010111101010) && ({row_reg, col_reg}<19'b1101100100100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1101100100100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1101100100100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1101100100100111010) && ({row_reg, col_reg}<19'b1101100100100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101100100100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1101100100100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101100100100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1101100100100111111) && ({row_reg, col_reg}<19'b1101100100101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101100100101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1101100100101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1101100100101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1101100100101010100) && ({row_reg, col_reg}<19'b1101100100111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1101100100111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1101100100111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1101100100111010000) && ({row_reg, col_reg}<19'b1101100100111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101100100111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1101100100111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1101100100111101010) && ({row_reg, col_reg}<19'b1101100110100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1101100110100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1101100110100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1101100110100111010) && ({row_reg, col_reg}<19'b1101100110100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101100110100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1101100110100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101100110100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1101100110100111111) && ({row_reg, col_reg}<19'b1101100110101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101100110101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1101100110101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1101100110101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1101100110101010100) && ({row_reg, col_reg}<19'b1101100110111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1101100110111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1101100110111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1101100110111010000) && ({row_reg, col_reg}<19'b1101100110111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101100110111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1101100110111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1101100110111101010) && ({row_reg, col_reg}<19'b1101101000100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1101101000100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1101101000100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1101101000100111010) && ({row_reg, col_reg}<19'b1101101000100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101101000100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1101101000100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101101000100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1101101000100111111) && ({row_reg, col_reg}<19'b1101101000101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101101000101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1101101000101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1101101000101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1101101000101010100) && ({row_reg, col_reg}<19'b1101101000111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1101101000111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1101101000111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1101101000111010000) && ({row_reg, col_reg}<19'b1101101000111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101101000111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1101101000111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1101101000111101010) && ({row_reg, col_reg}<19'b1101101010100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1101101010100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1101101010100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1101101010100111010) && ({row_reg, col_reg}<19'b1101101010100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101101010100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1101101010100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101101010100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1101101010100111111) && ({row_reg, col_reg}<19'b1101101010101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101101010101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1101101010101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1101101010101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1101101010101010100) && ({row_reg, col_reg}<19'b1101101010111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1101101010111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1101101010111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1101101010111010000) && ({row_reg, col_reg}<19'b1101101010111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101101010111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1101101010111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1101101010111101010) && ({row_reg, col_reg}<19'b1101101100100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1101101100100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1101101100100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1101101100100111010) && ({row_reg, col_reg}<19'b1101101100100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101101100100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1101101100100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101101100100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1101101100100111111) && ({row_reg, col_reg}<19'b1101101100101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101101100101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1101101100101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1101101100101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1101101100101010100) && ({row_reg, col_reg}<19'b1101101100111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1101101100111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1101101100111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1101101100111010000) && ({row_reg, col_reg}<19'b1101101100111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101101100111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1101101100111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1101101100111101010) && ({row_reg, col_reg}<19'b1101101110100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1101101110100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1101101110100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1101101110100111010) && ({row_reg, col_reg}<19'b1101101110100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101101110100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1101101110100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101101110100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1101101110100111111) && ({row_reg, col_reg}<19'b1101101110101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101101110101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1101101110101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1101101110101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1101101110101010100) && ({row_reg, col_reg}<19'b1101101110111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1101101110111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1101101110111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1101101110111010000) && ({row_reg, col_reg}<19'b1101101110111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101101110111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1101101110111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1101101110111101010) && ({row_reg, col_reg}<19'b1101110000100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1101110000100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1101110000100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1101110000100111010) && ({row_reg, col_reg}<19'b1101110000100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101110000100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1101110000100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101110000100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1101110000100111111) && ({row_reg, col_reg}<19'b1101110000101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101110000101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1101110000101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1101110000101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1101110000101010100) && ({row_reg, col_reg}<19'b1101110000111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1101110000111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1101110000111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1101110000111010000) && ({row_reg, col_reg}<19'b1101110000111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101110000111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1101110000111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1101110000111101010) && ({row_reg, col_reg}<19'b1101110010100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1101110010100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1101110010100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1101110010100111010) && ({row_reg, col_reg}<19'b1101110010100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101110010100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1101110010100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101110010100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1101110010100111111) && ({row_reg, col_reg}<19'b1101110010101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101110010101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1101110010101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1101110010101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1101110010101010100) && ({row_reg, col_reg}<19'b1101110010111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1101110010111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1101110010111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1101110010111010000) && ({row_reg, col_reg}<19'b1101110010111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101110010111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1101110010111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1101110010111101010) && ({row_reg, col_reg}<19'b1101110100100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1101110100100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1101110100100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1101110100100111010) && ({row_reg, col_reg}<19'b1101110100100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101110100100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1101110100100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101110100100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1101110100100111111) && ({row_reg, col_reg}<19'b1101110100101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101110100101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1101110100101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1101110100101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1101110100101010100) && ({row_reg, col_reg}<19'b1101110100111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1101110100111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1101110100111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1101110100111010000) && ({row_reg, col_reg}<19'b1101110100111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101110100111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1101110100111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1101110100111101010) && ({row_reg, col_reg}<19'b1101110110100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1101110110100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1101110110100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1101110110100111010) && ({row_reg, col_reg}<19'b1101110110100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101110110100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1101110110100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101110110100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1101110110100111111) && ({row_reg, col_reg}<19'b1101110110101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101110110101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1101110110101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1101110110101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1101110110101010100) && ({row_reg, col_reg}<19'b1101110110111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1101110110111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1101110110111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1101110110111010000) && ({row_reg, col_reg}<19'b1101110110111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101110110111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1101110110111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1101110110111101010) && ({row_reg, col_reg}<19'b1101111000100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1101111000100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1101111000100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1101111000100111010) && ({row_reg, col_reg}<19'b1101111000100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101111000100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1101111000100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101111000100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1101111000100111111) && ({row_reg, col_reg}<19'b1101111000101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101111000101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1101111000101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1101111000101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1101111000101010100) && ({row_reg, col_reg}<19'b1101111000111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1101111000111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1101111000111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1101111000111010000) && ({row_reg, col_reg}<19'b1101111000111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101111000111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1101111000111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1101111000111101010) && ({row_reg, col_reg}<19'b1101111010100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1101111010100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1101111010100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1101111010100111010) && ({row_reg, col_reg}<19'b1101111010100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101111010100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1101111010100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101111010100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1101111010100111111) && ({row_reg, col_reg}<19'b1101111010101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101111010101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1101111010101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1101111010101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1101111010101010100) && ({row_reg, col_reg}<19'b1101111010111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1101111010111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1101111010111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1101111010111010000) && ({row_reg, col_reg}<19'b1101111010111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101111010111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1101111010111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1101111010111101010) && ({row_reg, col_reg}<19'b1101111100100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1101111100100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1101111100100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1101111100100111010) && ({row_reg, col_reg}<19'b1101111100100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101111100100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1101111100100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101111100100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1101111100100111111) && ({row_reg, col_reg}<19'b1101111100101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101111100101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1101111100101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1101111100101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1101111100101010100) && ({row_reg, col_reg}<19'b1101111100111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1101111100111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1101111100111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1101111100111010000) && ({row_reg, col_reg}<19'b1101111100111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101111100111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1101111100111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1101111100111101010) && ({row_reg, col_reg}<19'b1101111110100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1101111110100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1101111110100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1101111110100111010) && ({row_reg, col_reg}<19'b1101111110100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101111110100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1101111110100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101111110100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1101111110100111111) && ({row_reg, col_reg}<19'b1101111110101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101111110101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1101111110101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1101111110101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1101111110101010100) && ({row_reg, col_reg}<19'b1101111110111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1101111110111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1101111110111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1101111110111010000) && ({row_reg, col_reg}<19'b1101111110111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1101111110111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1101111110111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1101111110111101010) && ({row_reg, col_reg}<19'b1110000000100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1110000000100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1110000000100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1110000000100111010) && ({row_reg, col_reg}<19'b1110000000100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110000000100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1110000000100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110000000100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1110000000100111111) && ({row_reg, col_reg}<19'b1110000000101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110000000101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1110000000101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1110000000101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1110000000101010100) && ({row_reg, col_reg}<19'b1110000000111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1110000000111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1110000000111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1110000000111010000) && ({row_reg, col_reg}<19'b1110000000111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110000000111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1110000000111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1110000000111101010) && ({row_reg, col_reg}<19'b1110000010100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1110000010100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1110000010100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1110000010100111010) && ({row_reg, col_reg}<19'b1110000010100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110000010100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1110000010100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110000010100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1110000010100111111) && ({row_reg, col_reg}<19'b1110000010101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110000010101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1110000010101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1110000010101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1110000010101010100) && ({row_reg, col_reg}<19'b1110000010111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1110000010111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1110000010111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1110000010111010000) && ({row_reg, col_reg}<19'b1110000010111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110000010111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1110000010111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1110000010111101010) && ({row_reg, col_reg}<19'b1110000100100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1110000100100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1110000100100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1110000100100111010) && ({row_reg, col_reg}<19'b1110000100100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110000100100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1110000100100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110000100100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1110000100100111111) && ({row_reg, col_reg}<19'b1110000100101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110000100101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1110000100101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1110000100101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1110000100101010100) && ({row_reg, col_reg}<19'b1110000100111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1110000100111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1110000100111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1110000100111010000) && ({row_reg, col_reg}<19'b1110000100111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110000100111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1110000100111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1110000100111101010) && ({row_reg, col_reg}<19'b1110000110100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1110000110100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1110000110100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1110000110100111010) && ({row_reg, col_reg}<19'b1110000110100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110000110100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1110000110100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110000110100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1110000110100111111) && ({row_reg, col_reg}<19'b1110000110101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110000110101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1110000110101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1110000110101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1110000110101010100) && ({row_reg, col_reg}<19'b1110000110111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1110000110111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1110000110111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1110000110111010000) && ({row_reg, col_reg}<19'b1110000110111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110000110111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1110000110111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1110000110111101010) && ({row_reg, col_reg}<19'b1110001000100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1110001000100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1110001000100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1110001000100111010) && ({row_reg, col_reg}<19'b1110001000100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110001000100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1110001000100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110001000100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1110001000100111111) && ({row_reg, col_reg}<19'b1110001000101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110001000101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1110001000101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1110001000101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1110001000101010100) && ({row_reg, col_reg}<19'b1110001000111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1110001000111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1110001000111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1110001000111010000) && ({row_reg, col_reg}<19'b1110001000111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110001000111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1110001000111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1110001000111101010) && ({row_reg, col_reg}<19'b1110001010100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1110001010100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1110001010100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1110001010100111010) && ({row_reg, col_reg}<19'b1110001010100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110001010100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1110001010100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110001010100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1110001010100111111) && ({row_reg, col_reg}<19'b1110001010101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110001010101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1110001010101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1110001010101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1110001010101010100) && ({row_reg, col_reg}<19'b1110001010111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1110001010111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1110001010111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1110001010111010000) && ({row_reg, col_reg}<19'b1110001010111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110001010111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1110001010111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1110001010111101010) && ({row_reg, col_reg}<19'b1110001100100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1110001100100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1110001100100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1110001100100111010) && ({row_reg, col_reg}<19'b1110001100100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110001100100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1110001100100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110001100100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1110001100100111111) && ({row_reg, col_reg}<19'b1110001100101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110001100101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1110001100101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1110001100101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1110001100101010100) && ({row_reg, col_reg}<19'b1110001100111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1110001100111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1110001100111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1110001100111010000) && ({row_reg, col_reg}<19'b1110001100111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110001100111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1110001100111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1110001100111101010) && ({row_reg, col_reg}<19'b1110001110100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1110001110100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1110001110100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1110001110100111010) && ({row_reg, col_reg}<19'b1110001110100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110001110100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1110001110100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110001110100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1110001110100111111) && ({row_reg, col_reg}<19'b1110001110101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110001110101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1110001110101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1110001110101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1110001110101010100) && ({row_reg, col_reg}<19'b1110001110111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1110001110111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1110001110111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1110001110111010000) && ({row_reg, col_reg}<19'b1110001110111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110001110111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1110001110111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1110001110111101010) && ({row_reg, col_reg}<19'b1110010000100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1110010000100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1110010000100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1110010000100111010) && ({row_reg, col_reg}<19'b1110010000100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110010000100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1110010000100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110010000100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1110010000100111111) && ({row_reg, col_reg}<19'b1110010000101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110010000101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1110010000101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1110010000101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1110010000101010100) && ({row_reg, col_reg}<19'b1110010000111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1110010000111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1110010000111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1110010000111010000) && ({row_reg, col_reg}<19'b1110010000111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110010000111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1110010000111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1110010000111101010) && ({row_reg, col_reg}<19'b1110010010100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1110010010100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1110010010100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1110010010100111010) && ({row_reg, col_reg}<19'b1110010010100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110010010100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1110010010100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110010010100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1110010010100111111) && ({row_reg, col_reg}<19'b1110010010101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110010010101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1110010010101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1110010010101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1110010010101010100) && ({row_reg, col_reg}<19'b1110010010111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1110010010111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1110010010111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1110010010111010000) && ({row_reg, col_reg}<19'b1110010010111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110010010111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1110010010111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1110010010111101010) && ({row_reg, col_reg}<19'b1110010100100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1110010100100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1110010100100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1110010100100111010) && ({row_reg, col_reg}<19'b1110010100100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110010100100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1110010100100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110010100100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1110010100100111111) && ({row_reg, col_reg}<19'b1110010100101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110010100101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1110010100101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1110010100101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1110010100101010100) && ({row_reg, col_reg}<19'b1110010100111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1110010100111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1110010100111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1110010100111010000) && ({row_reg, col_reg}<19'b1110010100111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110010100111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1110010100111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1110010100111101010) && ({row_reg, col_reg}<19'b1110010110100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1110010110100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1110010110100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1110010110100111010) && ({row_reg, col_reg}<19'b1110010110100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110010110100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1110010110100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110010110100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1110010110100111111) && ({row_reg, col_reg}<19'b1110010110101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110010110101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1110010110101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1110010110101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1110010110101010100) && ({row_reg, col_reg}<19'b1110010110111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1110010110111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1110010110111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1110010110111010000) && ({row_reg, col_reg}<19'b1110010110111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110010110111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1110010110111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1110010110111101010) && ({row_reg, col_reg}<19'b1110011000100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1110011000100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1110011000100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1110011000100111010) && ({row_reg, col_reg}<19'b1110011000100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110011000100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1110011000100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110011000100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1110011000100111111) && ({row_reg, col_reg}<19'b1110011000101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110011000101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1110011000101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1110011000101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1110011000101010100) && ({row_reg, col_reg}<19'b1110011000111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1110011000111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1110011000111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1110011000111010000) && ({row_reg, col_reg}<19'b1110011000111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110011000111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1110011000111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1110011000111101010) && ({row_reg, col_reg}<19'b1110011010100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1110011010100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1110011010100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1110011010100111010) && ({row_reg, col_reg}<19'b1110011010100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110011010100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1110011010100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110011010100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1110011010100111111) && ({row_reg, col_reg}<19'b1110011010101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110011010101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1110011010101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1110011010101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1110011010101010100) && ({row_reg, col_reg}<19'b1110011010111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1110011010111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1110011010111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1110011010111010000) && ({row_reg, col_reg}<19'b1110011010111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110011010111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1110011010111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1110011010111101010) && ({row_reg, col_reg}<19'b1110011100100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1110011100100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1110011100100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1110011100100111010) && ({row_reg, col_reg}<19'b1110011100100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110011100100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1110011100100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110011100100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1110011100100111111) && ({row_reg, col_reg}<19'b1110011100101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110011100101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1110011100101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1110011100101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1110011100101010100) && ({row_reg, col_reg}<19'b1110011100111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1110011100111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1110011100111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1110011100111010000) && ({row_reg, col_reg}<19'b1110011100111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110011100111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1110011100111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1110011100111101010) && ({row_reg, col_reg}<19'b1110011110100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1110011110100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1110011110100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1110011110100111010) && ({row_reg, col_reg}<19'b1110011110100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110011110100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1110011110100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110011110100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1110011110100111111) && ({row_reg, col_reg}<19'b1110011110101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110011110101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1110011110101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1110011110101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1110011110101010100) && ({row_reg, col_reg}<19'b1110011110111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1110011110111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1110011110111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1110011110111010000) && ({row_reg, col_reg}<19'b1110011110111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110011110111101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1110011110111101001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1110011110111101010) && ({row_reg, col_reg}<19'b1110100000100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1110100000100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1110100000100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1110100000100111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110100000100111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1110100000100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b1110100000100111101) && ({row_reg, col_reg}<19'b1110100000101000000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1110100000101000000) && ({row_reg, col_reg}<19'b1110100000101010000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b1110100000101010000) && ({row_reg, col_reg}<19'b1110100000101010010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1110100000101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1110100000101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1110100000101010100) && ({row_reg, col_reg}<19'b1110100000111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1110100000111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1110100000111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1110100000111010000) && ({row_reg, col_reg}<19'b1110100000111100000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110100000111100000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1110100000111100001) && ({row_reg, col_reg}<19'b1110100000111100011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b1110100000111100011) && ({row_reg, col_reg}<19'b1110100000111100101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1110100000111100101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110100000111100110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1110100000111100111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110100000111101000)) color_data = 12'b101010101010;

		if(({row_reg, col_reg}>=19'b1110100000111101001) && ({row_reg, col_reg}<19'b1110100010100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1110100010100111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1110100010100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1110100010100111010) && ({row_reg, col_reg}<19'b1110100010101010010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110100010101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1110100010101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1110100010101010100) && ({row_reg, col_reg}<19'b1110100010111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1110100010111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1110100010111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1110100010111010000) && ({row_reg, col_reg}<19'b1110100010111100000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110100010111100000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1110100010111100001) && ({row_reg, col_reg}<19'b1110100010111101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110100010111101000)) color_data = 12'b101010101010;

		if(({row_reg, col_reg}>=19'b1110100010111101001) && ({row_reg, col_reg}<19'b1110100100100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1110100100100111000)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1110100100100111001) && ({row_reg, col_reg}<19'b1110100100100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1110100100100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110100100100111101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1110100100100111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110100100100111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1110100100101000000) && ({row_reg, col_reg}<19'b1110100100101010010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110100100101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1110100100101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1110100100101010100) && ({row_reg, col_reg}<19'b1110100100111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1110100100111001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1110100100111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1110100100111010000) && ({row_reg, col_reg}<19'b1110100100111100010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110100100111100010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1110100100111100011) && ({row_reg, col_reg}<19'b1110100100111100111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110100100111100111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1110100100111101000)) color_data = 12'b101010101010;

		if(({row_reg, col_reg}>=19'b1110100100111101001) && ({row_reg, col_reg}<19'b1110100110100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1110100110100111000)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1110100110100111001) && ({row_reg, col_reg}<19'b1110100110100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1110100110100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110100110100111101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1110100110100111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110100110100111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1110100110101000000) && ({row_reg, col_reg}<19'b1110100110101010000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b1110100110101010000) && ({row_reg, col_reg}<19'b1110100110101010010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1110100110101010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1110100110101010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1110100110101010100) && ({row_reg, col_reg}<19'b1110100110111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1110100110111001110)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1110100110111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1110100110111010000) && ({row_reg, col_reg}<19'b1110100110111100010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110100110111100010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1110100110111100011) && ({row_reg, col_reg}<19'b1110100110111100101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110100110111100101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1110100110111100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110100110111100111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1110100110111101000)) color_data = 12'b101010101010;

		if(({row_reg, col_reg}>=19'b1110100110111101001) && ({row_reg, col_reg}<19'b1110101000100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1110101000100111000)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b1110101000100111001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1110101000100111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110101000100111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1110101000100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110101000100111101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1110101000100111110) && ({row_reg, col_reg}<19'b1110101000101010000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b1110101000101010000) && ({row_reg, col_reg}<19'b1110101000101010010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1110101000101010010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1110101000101010011)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=19'b1110101000101010100) && ({row_reg, col_reg}<19'b1110101000111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1110101000111001110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b1110101000111001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1110101000111010000) && ({row_reg, col_reg}<19'b1110101000111100010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110101000111100010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1110101000111100011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b1110101000111100100) && ({row_reg, col_reg}<19'b1110101000111100110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1110101000111100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110101000111100111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1110101000111101000)) color_data = 12'b101110111011;

		if(({row_reg, col_reg}>=19'b1110101000111101001) && ({row_reg, col_reg}<19'b1110101010100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1110101010100111000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b1110101010100111001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=19'b1110101010100111010) && ({row_reg, col_reg}<19'b1110101010100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1110101010100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110101010100111101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1110101010100111110) && ({row_reg, col_reg}<19'b1110101010101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110101010101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1110101010101010010)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=19'b1110101010101010011) && ({row_reg, col_reg}<19'b1110101010111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1110101010111001110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b1110101010111001111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=19'b1110101010111010000) && ({row_reg, col_reg}<19'b1110101010111100000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110101010111100000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1110101010111100001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110101010111100010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1110101010111100011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b1110101010111100100) && ({row_reg, col_reg}<19'b1110101010111100110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1110101010111100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110101010111100111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1110101010111101000)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=19'b1110101010111101001) && ({row_reg, col_reg}<19'b1110101100100111001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1110101100100111001)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=19'b1110101100100111010) && ({row_reg, col_reg}<19'b1110101100101000000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1110101100101000000) && ({row_reg, col_reg}<19'b1110101100101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110101100101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1110101100101010010)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=19'b1110101100101010011) && ({row_reg, col_reg}<19'b1110101100111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1110101100111001110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b1110101100111001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=19'b1110101100111010000) && ({row_reg, col_reg}<19'b1110101100111010011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1110101100111010011) && ({row_reg, col_reg}<19'b1110101100111100000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110101100111100000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1110101100111100001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110101100111100010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1110101100111100011) && ({row_reg, col_reg}<19'b1110101100111100111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110101100111100111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1110101100111101000)) color_data = 12'b110111011101;

		if(({row_reg, col_reg}>=19'b1110101100111101001) && ({row_reg, col_reg}<19'b1110101110100111001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1110101110100111001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1110101110100111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1110101110100111011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110101110100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1110101110100111101) && ({row_reg, col_reg}<19'b1110101110101010000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110101110101010000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1110101110101010001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1110101110101010010)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1110101110101010011) && ({row_reg, col_reg}<19'b1110101110111001111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1110101110111001111)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=19'b1110101110111010000) && ({row_reg, col_reg}<19'b1110101110111010011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1110101110111010011) && ({row_reg, col_reg}<19'b1110101110111100010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110101110111100010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1110101110111100011) && ({row_reg, col_reg}<19'b1110101110111100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110101110111100110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1110101110111100111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1110101110111101000)) color_data = 12'b110111011101;

		if(({row_reg, col_reg}>=19'b1110101110111101001) && ({row_reg, col_reg}<19'b1110110000100111001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1110110000100111001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b1110110000100111010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=19'b1110110000100111011) && ({row_reg, col_reg}<19'b1110110000100111101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1110110000100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110110000100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1110110000100111111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110110000101000000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1110110000101000001) && ({row_reg, col_reg}<19'b1110110000101000100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b1110110000101000100) && ({row_reg, col_reg}<19'b1110110000101000111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1110110000101000111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110110000101001000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1110110000101001001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110110000101001010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1110110000101001011) && ({row_reg, col_reg}<19'b1110110000101001110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110110000101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1110110000101001111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110110000101010000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1110110000101010001)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1110110000101010010)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=19'b1110110000101010011) && ({row_reg, col_reg}<19'b1110110000111001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1110110000111001110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b1110110000111001111)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b1110110000111010000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1110110000111010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b1110110000111010010) && ({row_reg, col_reg}<19'b1110110000111010100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1110110000111010100) && ({row_reg, col_reg}<19'b1110110000111010110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110110000111010110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1110110000111010111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b1110110000111011000) && ({row_reg, col_reg}<19'b1110110000111011010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1110110000111011010) && ({row_reg, col_reg}<19'b1110110000111011111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b1110110000111011111) && ({row_reg, col_reg}<19'b1110110000111100001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1110110000111100001) && ({row_reg, col_reg}<19'b1110110000111100100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110110000111100100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1110110000111100101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110110000111100110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1110110000111100111)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=19'b1110110000111101000) && ({row_reg, col_reg}<19'b1110110010100111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1110110010100111000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b1110110010100111001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1110110010100111010)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1110110010100111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1110110010100111100) && ({row_reg, col_reg}<19'b1110110010101000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b1110110010101000001) && ({row_reg, col_reg}<19'b1110110010101000011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1110110010101000011) && ({row_reg, col_reg}<19'b1110110010101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b1110110010101001100) && ({row_reg, col_reg}<19'b1110110010101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1110110010101001110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110110010101001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1110110010101010000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1110110010101010001)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1110110010101010010) && ({row_reg, col_reg}<19'b1110110010111001111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1110110010111001111)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b1110110010111010000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1110110010111010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1110110010111010010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b1110110010111010011) && ({row_reg, col_reg}<19'b1110110010111010101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1110110010111010101) && ({row_reg, col_reg}<19'b1110110010111010111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110110010111010111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1110110010111011000) && ({row_reg, col_reg}<19'b1110110010111011011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b1110110010111011011) && ({row_reg, col_reg}<19'b1110110010111011110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1110110010111011110) && ({row_reg, col_reg}<19'b1110110010111100000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b1110110010111100000) && ({row_reg, col_reg}<19'b1110110010111100110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1110110010111100110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1110110010111100111)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1110110010111101000) && ({row_reg, col_reg}<19'b1110110100100111010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1110110100100111010)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b1110110100100111011)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=19'b1110110100100111100) && ({row_reg, col_reg}<19'b1110110100101000010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1110110100101000010) && ({row_reg, col_reg}<19'b1110110100101000100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b1110110100101000100) && ({row_reg, col_reg}<19'b1110110100101001000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1110110100101001000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b1110110100101001001) && ({row_reg, col_reg}<19'b1110110100101001011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1110110100101001011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b1110110100101001100) && ({row_reg, col_reg}<19'b1110110100101010000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1110110100101010000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1110110100101010001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=19'b1110110100101010010) && ({row_reg, col_reg}<19'b1110110100111010000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1110110100111010000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b1110110100111010001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=19'b1110110100111010010) && ({row_reg, col_reg}<19'b1110110100111010100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110110100111010100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1110110100111010101) && ({row_reg, col_reg}<19'b1110110100111010111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b1110110100111010111) && ({row_reg, col_reg}<19'b1110110100111011001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1110110100111011001) && ({row_reg, col_reg}<19'b1110110100111011111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110110100111011111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1110110100111100000) && ({row_reg, col_reg}<19'b1110110100111100011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110110100111100011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1110110100111100100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110110100111100101)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1110110100111100110)) color_data = 12'b110111011101;

		if(({row_reg, col_reg}>=19'b1110110100111100111) && ({row_reg, col_reg}<19'b1110110110100111011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1110110110100111011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b1110110110100111100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1110110110100111101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1110110110100111110) && ({row_reg, col_reg}<19'b1110110110101001011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b1110110110101001011) && ({row_reg, col_reg}<19'b1110110110101001101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1110110110101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110110110101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1110110110101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1110110110101010000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=19'b1110110110101010001) && ({row_reg, col_reg}<19'b1110110110111010001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1110110110111010001)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b1110110110111010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=19'b1110110110111010011) && ({row_reg, col_reg}<19'b1110110110111010110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110110110111010110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1110110110111010111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b1110110110111011000) && ({row_reg, col_reg}<19'b1110110110111011110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1110110110111011110) && ({row_reg, col_reg}<19'b1110110110111100001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110110110111100001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1110110110111100010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b1110110110111100011) && ({row_reg, col_reg}<19'b1110110110111100101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1110110110111100101)) color_data = 12'b101110111011;

		if(({row_reg, col_reg}>=19'b1110110110111100110) && ({row_reg, col_reg}<19'b1110111000100111100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1110111000100111100)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b1110111000100111101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1110111000100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1110111000100111111) && ({row_reg, col_reg}<19'b1110111000101000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b1110111000101000001) && ({row_reg, col_reg}<19'b1110111000101000100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1110111000101000100) && ({row_reg, col_reg}<19'b1110111000101000111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b1110111000101000111) && ({row_reg, col_reg}<19'b1110111000101001001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1110111000101001001) && ({row_reg, col_reg}<19'b1110111000101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110111000101001101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1110111000101001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1110111000101001111)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=19'b1110111000101010000) && ({row_reg, col_reg}<19'b1110111000111010010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1110111000111010010)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1110111000111010011)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1110111000111010100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1110111000111010101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b1110111000111010110) && ({row_reg, col_reg}<19'b1110111000111011000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1110111000111011000) && ({row_reg, col_reg}<19'b1110111000111100000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110111000111100000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1110111000111100001) && ({row_reg, col_reg}<19'b1110111000111100011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110111000111100011)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1110111000111100100)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1110111000111100101)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1110111000111100110) && ({row_reg, col_reg}<19'b1110111010100111010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1110111010100111010)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=19'b1110111010100111011) && ({row_reg, col_reg}<19'b1110111010100111101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1110111010100111101)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b1110111010100111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1110111010100111111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1110111010101000000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1110111010101000001) && ({row_reg, col_reg}<19'b1110111010101000100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110111010101000100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1110111010101000101) && ({row_reg, col_reg}<19'b1110111010101000111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110111010101000111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1110111010101001000) && ({row_reg, col_reg}<19'b1110111010101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==19'b1110111010101001100)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1110111010101001101)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=19'b1110111010101001110) && ({row_reg, col_reg}<19'b1110111010111010011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1110111010111010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b1110111010111010100)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1110111010111010101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1110111010111010110) && ({row_reg, col_reg}<19'b1110111010111011011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b1110111010111011011) && ({row_reg, col_reg}<19'b1110111010111100010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1110111010111100010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1110111010111100011)) color_data = 12'b110111011101;

		if(({row_reg, col_reg}>=19'b1110111010111100100) && ({row_reg, col_reg}<19'b1110111100100111111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1110111100100111111)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1110111100101000000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1110111100101000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=19'b1110111100101000010) && ({row_reg, col_reg}<19'b1110111100101000101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=19'b1110111100101000101) && ({row_reg, col_reg}<19'b1110111100101000111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b1110111100101000111) && ({row_reg, col_reg}<19'b1110111100101001010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1110111100101001010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1110111100101001011)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1110111100101001100)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=19'b1110111100101001101) && ({row_reg, col_reg}<19'b1110111100111010100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1110111100111010100)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b1110111100111010101)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1110111100111010110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=19'b1110111100111010111) && ({row_reg, col_reg}<19'b1110111100111011011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1110111100111011011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=19'b1110111100111011100) && ({row_reg, col_reg}<19'b1110111100111100000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1110111100111100000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1110111100111100001)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1110111100111100010)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1110111100111100011) && ({row_reg, col_reg}<19'b1110111110101000000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1110111110101000000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b1110111110101000001)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b1110111110101000010)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1110111110101000011)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1110111110101000100)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=19'b1110111110101000101) && ({row_reg, col_reg}<19'b1110111110101000111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1110111110101000111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==19'b1110111110101001000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1110111110101001001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1110111110101001010)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b1110111110101001011)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=19'b1110111110101001100) && ({row_reg, col_reg}<19'b1110111110111010110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==19'b1110111110111010110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==19'b1110111110111010111)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1110111110111011000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1110111110111011001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1110111110111011010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=19'b1110111110111011011) && ({row_reg, col_reg}<19'b1110111110111011101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==19'b1110111110111011101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==19'b1110111110111011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==19'b1110111110111011111)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==19'b1110111110111100000)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==19'b1110111110111100001)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=19'b1110111110111100010) && ({row_reg, col_reg}<=19'b1110111111001111111)) color_data = 12'b111111111111;
	end
endmodule