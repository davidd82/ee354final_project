module tictactoeboard_rom
	(
		input wire clk,
		input wire [9:0] row,
		input wire [9:0] col,
		output reg [11:0] color_data
	);

	(* rom_style = "block" *)

	//signal declaration
	reg [9:0] row_reg;
	reg [9:0] col_reg;

	always @(posedge clk)
		begin
		row_reg <= row;
		col_reg <= col;
		end

	always @(*) begin
		if(({row_reg, col_reg}>=20'b00000000000000000000) && ({row_reg, col_reg}<20'b00000000000100101110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00000000000100101110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=20'b00000000000100101111) && ({row_reg, col_reg}<20'b00000000000100110001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00000000000100110001)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00000000000100110010)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==20'b00000000000100110011)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00000000000100110100)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=20'b00000000000100110101) && ({row_reg, col_reg}<20'b00000000000100111000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00000000000100111000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==20'b00000000000100111001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==20'b00000000000100111010)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00000000000100111011)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=20'b00000000000100111100) && ({row_reg, col_reg}<20'b00000000000100111110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00000000000100111110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00000000000100111111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=20'b00000000000101000000) && ({row_reg, col_reg}<20'b00000000000101000011)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=20'b00000000000101000011) && ({row_reg, col_reg}<20'b00000000000101000101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=20'b00000000000101000101) && ({row_reg, col_reg}<20'b00000000000101001001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00000000000101001001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=20'b00000000000101001010) && ({row_reg, col_reg}<20'b00000000001001000110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=20'b00000000001001000110) && ({row_reg, col_reg}<20'b00000000001001001000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=20'b00000000001001001000) && ({row_reg, col_reg}<20'b00000000001001001010)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00000000001001001010)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00000000001001001011)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00000000001001001100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==20'b00000000001001001101)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=20'b00000000001001001110) && ({row_reg, col_reg}<20'b00000000001001010000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00000000001001010000) && ({row_reg, col_reg}<20'b00000000001001010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==20'b00000000001001010010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==20'b00000000001001010011)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00000000001001010100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==20'b00000000001001010101)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=20'b00000000001001010110) && ({row_reg, col_reg}<20'b00000000001001100010)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=20'b00000000001001100010) && ({row_reg, col_reg}<20'b00000000001001100100)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00000000001001100100) && ({row_reg, col_reg}<20'b00000000010100100001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=20'b00000000010100100001) && ({row_reg, col_reg}<20'b00000000010100100011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=20'b00000000010100100011) && ({row_reg, col_reg}<20'b00000000010100100111)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00000000010100100111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=20'b00000000010100101000) && ({row_reg, col_reg}<20'b00000000010100101101)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00000000010100101101)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00000000010100101110)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=20'b00000000010100101111) && ({row_reg, col_reg}<20'b00000000010100110001)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00000000010100110001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00000000010100110010) && ({row_reg, col_reg}<20'b00000000010100110100)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=20'b00000000010100110100) && ({row_reg, col_reg}<20'b00000000010100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00000000010100111001) && ({row_reg, col_reg}<20'b00000000010100111011)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=20'b00000000010100111011) && ({row_reg, col_reg}<20'b00000000010100111110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00000000010100111110) && ({row_reg, col_reg}<20'b00000000010101000000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00000000010101000000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==20'b00000000010101000001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00000000010101000010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=20'b00000000010101000011) && ({row_reg, col_reg}<20'b00000000010101000101)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=20'b00000000010101000101) && ({row_reg, col_reg}<20'b00000000010101001000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=20'b00000000010101001000) && ({row_reg, col_reg}<20'b00000000011000111000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00000000011000111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=20'b00000000011000111001) && ({row_reg, col_reg}<20'b00000000011001000010)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=20'b00000000011001000010) && ({row_reg, col_reg}<20'b00000000011001000100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==20'b00000000011001000100)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00000000011001000101)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=20'b00000000011001000110) && ({row_reg, col_reg}<20'b00000000011001001000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=20'b00000000011001001000) && ({row_reg, col_reg}<20'b00000000011001001010)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00000000011001001010) && ({row_reg, col_reg}<20'b00000000011001001100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==20'b00000000011001001100)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=20'b00000000011001001101) && ({row_reg, col_reg}<20'b00000000011001010010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00000000011001010010) && ({row_reg, col_reg}<20'b00000000011001010100)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=20'b00000000011001010100) && ({row_reg, col_reg}<20'b00000000011001010110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00000000011001010110) && ({row_reg, col_reg}<20'b00000000011001011000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00000000011001011000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==20'b00000000011001011001)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=20'b00000000011001011010) && ({row_reg, col_reg}<20'b00000000011001011100)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00000000011001011100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=20'b00000000011001011101) && ({row_reg, col_reg}<20'b00000000011001011111)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00000000011001011111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=20'b00000000011001100000) && ({row_reg, col_reg}<20'b00000000011001100111)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00000000011001100111)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00000000011001101000) && ({row_reg, col_reg}<20'b00000000100100100100)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00000000100100100100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=20'b00000000100100100101) && ({row_reg, col_reg}<20'b00000000100100101011)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00000000100100101011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00000000100100101100)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00000000100100101101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==20'b00000000100100101110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=20'b00000000100100101111) && ({row_reg, col_reg}<20'b00000000100100110100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00000000100100110100) && ({row_reg, col_reg}<20'b00000000100100111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00000000100100111110) && ({row_reg, col_reg}<20'b00000000100101000000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00000000100101000000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==20'b00000000100101000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==20'b00000000100101000010)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00000000100101000011)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=20'b00000000100101000100) && ({row_reg, col_reg}<20'b00000000100101000110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=20'b00000000100101000110) && ({row_reg, col_reg}<20'b00000000100101001000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00000000100101001000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=20'b00000000100101001001) && ({row_reg, col_reg}<20'b00000000100101001011)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00000000100101001011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=20'b00000000100101001100) && ({row_reg, col_reg}<20'b00000000101001000000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00000000101001000000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=20'b00000000101001000001) && ({row_reg, col_reg}<20'b00000000101001000100)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00000000101001000100)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00000000101001000101)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00000000101001000110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00000000101001000111) && ({row_reg, col_reg}<20'b00000000101001001010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00000000101001001010) && ({row_reg, col_reg}<20'b00000000101001010110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00000000101001010110) && ({row_reg, col_reg}<20'b00000000101001011001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00000000101001011001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==20'b00000000101001011010)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==20'b00000000101001011011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=20'b00000000101001011100) && ({row_reg, col_reg}<20'b00000000101001100111)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00000000101001100111)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00000000101001101000) && ({row_reg, col_reg}<20'b00000000110100100000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00000000110100100000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=20'b00000000110100100001) && ({row_reg, col_reg}<20'b00000000110100100011)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=20'b00000000110100100011) && ({row_reg, col_reg}<20'b00000000110100100101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=20'b00000000110100100101) && ({row_reg, col_reg}<20'b00000000110100101010)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00000000110100101010)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==20'b00000000110100101011)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00000000110100101100) && ({row_reg, col_reg}<20'b00000000110100101111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00000000110100101111) && ({row_reg, col_reg}<20'b00000000110100110101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00000000110100110101) && ({row_reg, col_reg}<20'b00000000110100110111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00000000110100110111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00000000110100111000) && ({row_reg, col_reg}<20'b00000000110100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00000000110100111100) && ({row_reg, col_reg}<20'b00000000110101000000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00000000110101000000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00000000110101000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==20'b00000000110101000010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==20'b00000000110101000011)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=20'b00000000110101000100) && ({row_reg, col_reg}<20'b00000000110101001011)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00000000110101001011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=20'b00000000110101001100) && ({row_reg, col_reg}<20'b00000000111001000011)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00000000111001000011)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==20'b00000000111001000100)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=20'b00000000111001000101) && ({row_reg, col_reg}<20'b00000000111001001001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00000000111001001001) && ({row_reg, col_reg}<20'b00000000111001001011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00000000111001001011) && ({row_reg, col_reg}<20'b00000000111001010100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00000000111001010100) && ({row_reg, col_reg}<20'b00000000111001011001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00000000111001011001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00000000111001011010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==20'b00000000111001011011)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00000000111001011100)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=20'b00000000111001011101) && ({row_reg, col_reg}<20'b00000000111001100100)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00000000111001100100)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00000000111001100101) && ({row_reg, col_reg}<20'b00000001000100101000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00000001000100101000)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00000001000100101001)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00000001000100101010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==20'b00000001000100101011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00000001000100101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00000001000100101101) && ({row_reg, col_reg}<20'b00000001000100101111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00000001000100101111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00000001000100110000) && ({row_reg, col_reg}<20'b00000001000100110100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00000001000100110100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00000001000100110101) && ({row_reg, col_reg}<20'b00000001000100110111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00000001000100110111) && ({row_reg, col_reg}<20'b00000001000100111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00000001000100111100) && ({row_reg, col_reg}<20'b00000001000100111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00000001000100111110) && ({row_reg, col_reg}<20'b00000001000101000010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00000001000101000010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00000001000101000011)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==20'b00000001000101000100)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00000001000101000101)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=20'b00000001000101000110) && ({row_reg, col_reg}<20'b00000001001001000001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00000001001001000001)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00000001001001000010)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00000001001001000011)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==20'b00000001001001000100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00000001001001000101) && ({row_reg, col_reg}<20'b00000001001001000111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00000001001001000111) && ({row_reg, col_reg}<20'b00000001001001001001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00000001001001001001) && ({row_reg, col_reg}<20'b00000001001001011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00000001001001011000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00000001001001011001) && ({row_reg, col_reg}<20'b00000001001001011011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00000001001001011011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00000001001001011100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==20'b00000001001001011101)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==20'b00000001001001011110)) color_data = 12'b110111011101;

		if(({row_reg, col_reg}>=20'b00000001001001011111) && ({row_reg, col_reg}<20'b00000001010100100001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=20'b00000001010100100001) && ({row_reg, col_reg}<20'b00000001010100100011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=20'b00000001010100100011) && ({row_reg, col_reg}<20'b00000001010100100101)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00000001010100100101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==20'b00000001010100100110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00000001010100100111)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==20'b00000001010100101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==20'b00000001010100101001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=20'b00000001010100101010) && ({row_reg, col_reg}<20'b00000001010100101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00000001010100101100) && ({row_reg, col_reg}<20'b00000001010100101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00000001010100101110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00000001010100101111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00000001010100110000) && ({row_reg, col_reg}<20'b00000001010100111000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00000001010100111000) && ({row_reg, col_reg}<20'b00000001010101000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00000001010101000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00000001010101000010) && ({row_reg, col_reg}<20'b00000001010101000101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00000001010101000101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00000001010101000110) && ({row_reg, col_reg}<20'b00000001010101001000)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00000001010101001000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=20'b00000001010101001001) && ({row_reg, col_reg}<20'b00000001010101001011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=20'b00000001010101001011) && ({row_reg, col_reg}<20'b00000001011000111101)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00000001011000111101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=20'b00000001011000111110) && ({row_reg, col_reg}<20'b00000001011001000000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00000001011001000000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==20'b00000001011001000001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00000001011001000010) && ({row_reg, col_reg}<20'b00000001011001000110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00000001011001000110) && ({row_reg, col_reg}<20'b00000001011001001000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00000001011001001000) && ({row_reg, col_reg}<20'b00000001011001001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00000001011001001111) && ({row_reg, col_reg}<20'b00000001011001010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00000001011001010001) && ({row_reg, col_reg}<20'b00000001011001010100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00000001011001010100) && ({row_reg, col_reg}<20'b00000001011001010110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00000001011001010110) && ({row_reg, col_reg}<20'b00000001011001011000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00000001011001011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00000001011001011001) && ({row_reg, col_reg}<20'b00000001011001011101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00000001011001011101)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==20'b00000001011001011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00000001011001011111)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=20'b00000001011001100000) && ({row_reg, col_reg}<20'b00000001011001100010)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00000001011001100010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00000001011001100011) && ({row_reg, col_reg}<20'b00000001100100100110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00000001100100100110)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==20'b00000001100100100111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==20'b00000001100100101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00000001100100101001) && ({row_reg, col_reg}<20'b00000001100100101011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00000001100100101011) && ({row_reg, col_reg}<20'b00000001100100101101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00000001100100101101) && ({row_reg, col_reg}<20'b00000001100100101111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00000001100100101111) && ({row_reg, col_reg}<20'b00000001100100110001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00000001100100110001) && ({row_reg, col_reg}<20'b00000001100100110011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00000001100100110011) && ({row_reg, col_reg}<20'b00000001100100111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00000001100100111010) && ({row_reg, col_reg}<20'b00000001100101000100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00000001100101000100) && ({row_reg, col_reg}<20'b00000001100101000110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00000001100101000110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==20'b00000001100101000111)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00000001100101001000)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00000001100101001001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00000001100101001010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=20'b00000001100101001011) && ({row_reg, col_reg}<20'b00000001101000111110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00000001101000111110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00000001101000111111)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==20'b00000001101001000000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=20'b00000001101001000001) && ({row_reg, col_reg}<20'b00000001101001000100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00000001101001000100) && ({row_reg, col_reg}<20'b00000001101001000111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00000001101001000111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00000001101001001000) && ({row_reg, col_reg}<20'b00000001101001001110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00000001101001001110) && ({row_reg, col_reg}<20'b00000001101001010000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00000001101001010000) && ({row_reg, col_reg}<20'b00000001101001011100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00000001101001011100) && ({row_reg, col_reg}<20'b00000001101001011111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00000001101001011111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==20'b00000001101001100000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==20'b00000001101001100001)) color_data = 12'b110111011101;

		if(({row_reg, col_reg}>=20'b00000001101001100010) && ({row_reg, col_reg}<20'b00000001110100100100)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00000001110100100100)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00000001110100100101)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00000001110100100110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==20'b00000001110100100111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00000001110100101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00000001110100101001) && ({row_reg, col_reg}<20'b00000001110100101011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00000001110100101011) && ({row_reg, col_reg}<20'b00000001110100101110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00000001110100101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00000001110100101111) && ({row_reg, col_reg}<20'b00000001110100110011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00000001110100110011) && ({row_reg, col_reg}<20'b00000001110100110101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00000001110100110101) && ({row_reg, col_reg}<20'b00000001110100111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00000001110100111010) && ({row_reg, col_reg}<20'b00000001110100111101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00000001110100111101) && ({row_reg, col_reg}<20'b00000001110101000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00000001110101000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00000001110101000010) && ({row_reg, col_reg}<20'b00000001110101000100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00000001110101000100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00000001110101000101) && ({row_reg, col_reg}<20'b00000001110101000111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00000001110101000111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==20'b00000001110101001000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00000001110101001001)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=20'b00000001110101001010) && ({row_reg, col_reg}<20'b00000001110101001100)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=20'b00000001110101001100) && ({row_reg, col_reg}<20'b00000001110101001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==20'b00000001110101001110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00000001110101001111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=20'b00000001110101010000) && ({row_reg, col_reg}<20'b00000001111000111101)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00000001111000111101)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00000001111000111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00000001111000111111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=20'b00000001111001000000) && ({row_reg, col_reg}<20'b00000001111001000010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00000001111001000010) && ({row_reg, col_reg}<20'b00000001111001000101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00000001111001000101) && ({row_reg, col_reg}<20'b00000001111001000111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00000001111001000111) && ({row_reg, col_reg}<20'b00000001111001001001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00000001111001001001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00000001111001001010) && ({row_reg, col_reg}<20'b00000001111001010101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00000001111001010101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00000001111001010110) && ({row_reg, col_reg}<20'b00000001111001011001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00000001111001011001) && ({row_reg, col_reg}<20'b00000001111001011011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00000001111001011011) && ({row_reg, col_reg}<20'b00000001111001011111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00000001111001011111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00000001111001100000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==20'b00000001111001100001)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=20'b00000001111001100010) && ({row_reg, col_reg}<20'b00000010000100100000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00000010000100100000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=20'b00000010000100100001) && ({row_reg, col_reg}<20'b00000010000100100100)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00000010000100100100)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00000010000100100101) && ({row_reg, col_reg}<20'b00000010000100100111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00000010000100100111) && ({row_reg, col_reg}<20'b00000010000101001000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00000010000101001000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==20'b00000010000101001001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=20'b00000010000101001010) && ({row_reg, col_reg}<20'b00000010000101001100)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00000010000101001100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=20'b00000010000101001101) && ({row_reg, col_reg}<20'b00000010000101001111)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00000010000101001111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=20'b00000010000101010000) && ({row_reg, col_reg}<20'b00000010001000111001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00000010001000111001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=20'b00000010001000111010) && ({row_reg, col_reg}<20'b00000010001000111101)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00000010001000111101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00000010001000111110) && ({row_reg, col_reg}<20'b00000010001001000000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00000010001001000000) && ({row_reg, col_reg}<20'b00000010001001100000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00000010001001100000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00000010001001100001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==20'b00000010001001100010)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=20'b00000010001001100011) && ({row_reg, col_reg}<20'b00000010010100100011)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00000010010100100011)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==20'b00000010010100100100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==20'b00000010010100100101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00000010010100100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00000010010100100111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00000010010100101000) && ({row_reg, col_reg}<20'b00000010010101001000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00000010010101001000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00000010010101001001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==20'b00000010010101001010)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00000010010101001011)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00000010010101001100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==20'b00000010010101001101)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00000010010101001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=20'b00000010010101001111) && ({row_reg, col_reg}<20'b00000010011000111010)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00000010011000111010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==20'b00000010011000111011)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00000010011000111100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==20'b00000010011000111101)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==20'b00000010011000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00000010011000111111) && ({row_reg, col_reg}<20'b00000010011001100000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00000010011001100000) && ({row_reg, col_reg}<20'b00000010011001100010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00000010011001100010)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00000010011001100011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=20'b00000010011001100100) && ({row_reg, col_reg}<20'b00000010011001100110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00000010011001100110)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00000010011001100111) && ({row_reg, col_reg}<20'b00000010100100100010)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00000010100100100010)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00000010100100100011)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00000010100100100100) && ({row_reg, col_reg}<20'b00000010100100100110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00000010100100100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00000010100100100111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00000010100100101000) && ({row_reg, col_reg}<20'b00000010100101001001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00000010100101001001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00000010100101001010)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00000010100101001011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=20'b00000010100101001100) && ({row_reg, col_reg}<20'b00000010100101001110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00000010100101001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=20'b00000010100101001111) && ({row_reg, col_reg}<20'b00000010101000111000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00000010101000111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==20'b00000010101000111001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00000010101000111010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==20'b00000010101000111011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00000010101000111100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==20'b00000010101000111101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00000010101000111110) && ({row_reg, col_reg}<20'b00000010101001100010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00000010101001100010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==20'b00000010101001100011)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00000010101001100100)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=20'b00000010101001100101) && ({row_reg, col_reg}<20'b00000010101001100111)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00000010101001100111) && ({row_reg, col_reg}<20'b00000010110100100010)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00000010110100100010)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==20'b00000010110100100011)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==20'b00000010110100100100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00000010110100100101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00000010110100100110) && ({row_reg, col_reg}<20'b00000010110101001000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00000010110101001000) && ({row_reg, col_reg}<20'b00000010110101001010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00000010110101001010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==20'b00000010110101001011)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=20'b00000010110101001100) && ({row_reg, col_reg}<20'b00000010110101001111)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00000010110101001111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=20'b00000010110101010000) && ({row_reg, col_reg}<20'b00000010111000111011)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00000010111000111011)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00000010111000111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00000010111000111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00000010111000111110) && ({row_reg, col_reg}<20'b00000010111001000000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00000010111001000000) && ({row_reg, col_reg}<20'b00000010111001100001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00000010111001100001) && ({row_reg, col_reg}<20'b00000010111001100011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00000010111001100011)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==20'b00000010111001100100)) color_data = 12'b110111011101;

		if(({row_reg, col_reg}>=20'b00000010111001100101) && ({row_reg, col_reg}<20'b00000011000100100001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00000011000100100001)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00000011000100100010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00000011000100100011) && ({row_reg, col_reg}<20'b00000011000100100101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00000011000100100101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00000011000100100110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00000011000100100111) && ({row_reg, col_reg}<20'b00000011000101001000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00000011000101001000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00000011000101001001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00000011000101001010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00000011000101001011)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==20'b00000011000101001100)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=20'b00000011000101001101) && ({row_reg, col_reg}<20'b00000011001000111010)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00000011001000111010)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==20'b00000011001000111011)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=20'b00000011001000111100) && ({row_reg, col_reg}<20'b00000011001000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00000011001000111110) && ({row_reg, col_reg}<20'b00000011001001100000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00000011001001100000) && ({row_reg, col_reg}<20'b00000011001001100010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00000011001001100010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00000011001001100011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00000011001001100100)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00000011001001100101)) color_data = 12'b110111011101;

		if(({row_reg, col_reg}>=20'b00000011001001100110) && ({row_reg, col_reg}<20'b00000011010100100001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00000011010100100001)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00000011010100100010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00000011010100100011) && ({row_reg, col_reg}<20'b00000011010100100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00000011010100100110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00000011010100100111) && ({row_reg, col_reg}<20'b00000011010101001000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00000011010101001000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00000011010101001001) && ({row_reg, col_reg}<20'b00000011010101001011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00000011010101001011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00000011010101001100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==20'b00000011010101001101)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00000011010101001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=20'b00000011010101001111) && ({row_reg, col_reg}<20'b00000011011000111000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00000011011000111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==20'b00000011011000111001)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00000011011000111010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==20'b00000011011000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00000011011000111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00000011011000111101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00000011011000111110) && ({row_reg, col_reg}<20'b00000011011001100000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00000011011001100000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00000011011001100001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00000011011001100010) && ({row_reg, col_reg}<20'b00000011011001100101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00000011011001100101)) color_data = 12'b101110111011;

		if(({row_reg, col_reg}>=20'b00000011011001100110) && ({row_reg, col_reg}<20'b00000011100100100000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00000011100100100000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==20'b00000011100100100001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==20'b00000011100100100010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00000011100100100011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00000011100100100100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00000011100100100101) && ({row_reg, col_reg}<20'b00000011100101001000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00000011100101001000) && ({row_reg, col_reg}<20'b00000011100101001010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00000011100101001010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00000011100101001011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00000011100101001100)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==20'b00000011100101001101)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=20'b00000011100101001110) && ({row_reg, col_reg}<20'b00000011101000111001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00000011101000111001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==20'b00000011101000111010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==20'b00000011101000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00000011101000111100) && ({row_reg, col_reg}<20'b00000011101000111111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00000011101000111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00000011101001000000) && ({row_reg, col_reg}<20'b00000011101001100000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00000011101001100000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00000011101001100001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00000011101001100010) && ({row_reg, col_reg}<20'b00000011101001100100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00000011101001100100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00000011101001100101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==20'b00000011101001100110)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=20'b00000011101001100111) && ({row_reg, col_reg}<20'b00000011110100100000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00000011110100100000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==20'b00000011110100100001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00000011110100100010) && ({row_reg, col_reg}<20'b00000011110100100100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00000011110100100100) && ({row_reg, col_reg}<20'b00000011110100100110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00000011110100100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00000011110100100111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00000011110100101000) && ({row_reg, col_reg}<20'b00000011110101001001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00000011110101001001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00000011110101001010) && ({row_reg, col_reg}<20'b00000011110101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00000011110101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00000011110101001101)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00000011110101001110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00000011110101001111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=20'b00000011110101010000) && ({row_reg, col_reg}<20'b00000011111000111000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00000011111000111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==20'b00000011111000111001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00000011111000111010) && ({row_reg, col_reg}<20'b00000011111000111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00000011111000111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00000011111000111101) && ({row_reg, col_reg}<20'b00000011111000111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00000011111000111111) && ({row_reg, col_reg}<20'b00000011111001100001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00000011111001100001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00000011111001100010) && ({row_reg, col_reg}<20'b00000011111001100101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00000011111001100101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00000011111001100110)) color_data = 12'b101110111011;

		if(({row_reg, col_reg}>=20'b00000011111001100111) && ({row_reg, col_reg}<20'b00000100000100011010)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00000100000100011010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=20'b00000100000100011011) && ({row_reg, col_reg}<20'b00000100000100011111)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00000100000100011111)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00000100000100100000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=20'b00000100000100100001) && ({row_reg, col_reg}<20'b00000100000100100100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00000100000100100100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00000100000100100101) && ({row_reg, col_reg}<20'b00000100000100100111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00000100000100100111) && ({row_reg, col_reg}<20'b00000100000101001000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00000100000101001000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00000100000101001001) && ({row_reg, col_reg}<20'b00000100000101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00000100000101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00000100000101001101)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==20'b00000100000101001110)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=20'b00000100000101001111) && ({row_reg, col_reg}<20'b00000100001000111000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00000100001000111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=20'b00000100001000111001) && ({row_reg, col_reg}<20'b00000100001000111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00000100001000111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00000100001000111101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00000100001000111110) && ({row_reg, col_reg}<20'b00000100001001100000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00000100001001100000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00000100001001100001) && ({row_reg, col_reg}<20'b00000100001001100011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00000100001001100011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00000100001001100100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00000100001001100101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00000100001001100110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==20'b00000100001001100111)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00000100001001101000)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00000100001001101001) && ({row_reg, col_reg}<20'b00000100010100011111)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00000100010100011111)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=20'b00000100010100100000) && ({row_reg, col_reg}<20'b00000100010100100010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00000100010100100010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00000100010100100011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00000100010100100100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00000100010100100101) && ({row_reg, col_reg}<20'b00000100010100100111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00000100010100100111) && ({row_reg, col_reg}<20'b00000100010101001000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00000100010101001000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00000100010101001001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00000100010101001010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00000100010101001011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00000100010101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00000100010101001101)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==20'b00000100010101001110)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=20'b00000100010101001111) && ({row_reg, col_reg}<20'b00000100011000111000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00000100011000111000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00000100011000111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00000100011000111010) && ({row_reg, col_reg}<20'b00000100011001100001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00000100011001100001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00000100011001100010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00000100011001100011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00000100011001100100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00000100011001100101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00000100011001100110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==20'b00000100011001100111)) color_data = 12'b110111011101;

		if(({row_reg, col_reg}>=20'b00000100011001101000) && ({row_reg, col_reg}<20'b00000100100100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00000100100100011110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00000100100100011111)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00000100100100100000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00000100100100100001) && ({row_reg, col_reg}<20'b00000100100100100101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00000100100100100101) && ({row_reg, col_reg}<20'b00000100100100100111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00000100100100100111) && ({row_reg, col_reg}<20'b00000100100101001010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00000100100101001010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00000100100101001011) && ({row_reg, col_reg}<20'b00000100100101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00000100100101001101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00000100100101001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00000100100101001111) && ({row_reg, col_reg}<20'b00000100101000111000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00000100101000111000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00000100101000111001) && ({row_reg, col_reg}<20'b00000100101000111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00000100101000111101) && ({row_reg, col_reg}<20'b00000100101000111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00000100101000111111) && ({row_reg, col_reg}<20'b00000100101001100001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00000100101001100001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00000100101001100010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00000100101001100011) && ({row_reg, col_reg}<20'b00000100101001100101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00000100101001100101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00000100101001100110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==20'b00000100101001100111)) color_data = 12'b110111011101;

		if(({row_reg, col_reg}>=20'b00000100101001101000) && ({row_reg, col_reg}<20'b00000100110100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00000100110100011110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00000100110100011111)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00000100110100100000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00000100110100100001) && ({row_reg, col_reg}<20'b00000100110100100101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00000100110100100101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00000100110100100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00000100110100100111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00000100110100101000) && ({row_reg, col_reg}<20'b00000100110101001010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00000100110101001010) && ({row_reg, col_reg}<20'b00000100110101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00000100110101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00000100110101001101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00000100110101001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00000100110101001111) && ({row_reg, col_reg}<20'b00000100111000110111)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00000100111000110111)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00000100111000111000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==20'b00000100111000111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00000100111000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00000100111000111011) && ({row_reg, col_reg}<20'b00000100111000111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00000100111000111111) && ({row_reg, col_reg}<20'b00000100111001100001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00000100111001100001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00000100111001100010) && ({row_reg, col_reg}<20'b00000100111001100100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00000100111001100100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00000100111001100101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00000100111001100110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00000100111001100111)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=20'b00000100111001101000) && ({row_reg, col_reg}<20'b00000101000100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00000101000100011110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00000101000100011111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00000101000100100000) && ({row_reg, col_reg}<20'b00000101000100100011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00000101000100100011) && ({row_reg, col_reg}<20'b00000101000100100101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00000101000100100101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00000101000100100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00000101000100100111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00000101000100101000) && ({row_reg, col_reg}<20'b00000101000101001000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00000101000101001000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00000101000101001001) && ({row_reg, col_reg}<20'b00000101000101001011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00000101000101001011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00000101000101001100) && ({row_reg, col_reg}<20'b00000101000101001110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00000101000101001110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00000101000101001111) && ({row_reg, col_reg}<20'b00000101001000110111)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00000101001000110111)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==20'b00000101001000111000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==20'b00000101001000111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00000101001000111010) && ({row_reg, col_reg}<20'b00000101001001100001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00000101001001100001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00000101001001100010) && ({row_reg, col_reg}<20'b00000101001001100100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00000101001001100100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00000101001001100101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00000101001001100110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00000101001001100111)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00000101001001101000)) color_data = 12'b110111011101;

		if(({row_reg, col_reg}>=20'b00000101001001101001) && ({row_reg, col_reg}<20'b00000101010100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00000101010100011110)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==20'b00000101010100011111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=20'b00000101010100100000) && ({row_reg, col_reg}<20'b00000101010100100011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00000101010100100011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00000101010100100100) && ({row_reg, col_reg}<20'b00000101010100100110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00000101010100100110) && ({row_reg, col_reg}<20'b00000101010101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00000101010101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00000101010101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00000101010101001110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==20'b00000101010101001111)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=20'b00000101010101010000) && ({row_reg, col_reg}<20'b00000101011000110001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00000101011000110001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=20'b00000101011000110010) && ({row_reg, col_reg}<20'b00000101011000110111)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00000101011000110111)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==20'b00000101011000111000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==20'b00000101011000111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00000101011000111010) && ({row_reg, col_reg}<20'b00000101011000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00000101011000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00000101011000111111) && ({row_reg, col_reg}<20'b00000101011001100101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00000101011001100101) && ({row_reg, col_reg}<20'b00000101011001100111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00000101011001100111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==20'b00000101011001101000)) color_data = 12'b110111011101;

		if(({row_reg, col_reg}>=20'b00000101011001101001) && ({row_reg, col_reg}<20'b00000101100100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00000101100100011110)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==20'b00000101100100011111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=20'b00000101100100100000) && ({row_reg, col_reg}<20'b00000101100100100011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00000101100100100011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00000101100100100100) && ({row_reg, col_reg}<20'b00000101100100100110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00000101100100100110) && ({row_reg, col_reg}<20'b00000101100101001001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00000101100101001001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00000101100101001010) && ({row_reg, col_reg}<20'b00000101100101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00000101100101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00000101100101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00000101100101001110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==20'b00000101100101001111)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=20'b00000101100101010000) && ({row_reg, col_reg}<20'b00000101101000110001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00000101101000110001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=20'b00000101101000110010) && ({row_reg, col_reg}<20'b00000101101000110111)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00000101101000110111)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00000101101000111000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=20'b00000101101000111001) && ({row_reg, col_reg}<20'b00000101101000111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00000101101000111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00000101101000111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00000101101000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00000101101000111111) && ({row_reg, col_reg}<20'b00000101101001100011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00000101101001100011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00000101101001100100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00000101101001100101) && ({row_reg, col_reg}<20'b00000101101001100111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00000101101001100111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==20'b00000101101001101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==20'b00000101101001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00000101101001101010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=20'b00000101101001101011) && ({row_reg, col_reg}<20'b00000101101001101110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00000101101001101110)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00000101101001101111) && ({row_reg, col_reg}<20'b00000101110100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00000101110100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00000101110100011111) && ({row_reg, col_reg}<20'b00000101110100100001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00000101110100100001) && ({row_reg, col_reg}<20'b00000101110100100100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00000101110100100100) && ({row_reg, col_reg}<20'b00000101110100100110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00000101110100100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00000101110100100111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00000101110100101000) && ({row_reg, col_reg}<20'b00000101110101001001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00000101110101001001) && ({row_reg, col_reg}<20'b00000101110101001011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00000101110101001011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00000101110101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00000101110101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00000101110101001110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==20'b00000101110101001111)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00000101110101010000) && ({row_reg, col_reg}<20'b00000101111000110001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00000101111000110001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=20'b00000101111000110010) && ({row_reg, col_reg}<20'b00000101111000110111)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00000101111000110111)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00000101111000111000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=20'b00000101111000111001) && ({row_reg, col_reg}<20'b00000101111000111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00000101111000111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00000101111000111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00000101111000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00000101111000111111) && ({row_reg, col_reg}<20'b00000101111001100000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00000101111001100000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00000101111001100001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00000101111001100010) && ({row_reg, col_reg}<20'b00000101111001100100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00000101111001100100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00000101111001100101) && ({row_reg, col_reg}<20'b00000101111001100111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00000101111001100111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==20'b00000101111001101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==20'b00000101111001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00000101111001101010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=20'b00000101111001101011) && ({row_reg, col_reg}<20'b00000101111001101110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00000101111001101110)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00000101111001101111) && ({row_reg, col_reg}<20'b00000110000100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00000110000100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00000110000100011111) && ({row_reg, col_reg}<20'b00000110000101001000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00000110000101001000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00000110000101001001) && ({row_reg, col_reg}<20'b00000110000101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00000110000101001100) && ({row_reg, col_reg}<20'b00000110000101001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00000110000101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00000110000101010000) && ({row_reg, col_reg}<20'b00000110001000110111)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00000110001000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00000110001000111000) && ({row_reg, col_reg}<20'b00000110001000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00000110001000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00000110001000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00000110001000111100) && ({row_reg, col_reg}<20'b00000110001000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00000110001000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00000110001000111111) && ({row_reg, col_reg}<20'b00000110001001100100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00000110001001100100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00000110001001100101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00000110001001100110) && ({row_reg, col_reg}<20'b00000110001001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00000110001001101000)) color_data = 12'b101110111011;

		if(({row_reg, col_reg}>=20'b00000110001001101001) && ({row_reg, col_reg}<20'b00000110010100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00000110010100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00000110010100011111) && ({row_reg, col_reg}<20'b00000110010101001000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00000110010101001000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00000110010101001001) && ({row_reg, col_reg}<20'b00000110010101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00000110010101001100) && ({row_reg, col_reg}<20'b00000110010101001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00000110010101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00000110010101010000) && ({row_reg, col_reg}<20'b00000110011000110111)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00000110011000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00000110011000111000) && ({row_reg, col_reg}<20'b00000110011000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00000110011000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00000110011000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00000110011000111100) && ({row_reg, col_reg}<20'b00000110011000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00000110011000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00000110011000111111) && ({row_reg, col_reg}<20'b00000110011001100100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00000110011001100100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00000110011001100101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00000110011001100110) && ({row_reg, col_reg}<20'b00000110011001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00000110011001101000)) color_data = 12'b101110111011;

		if(({row_reg, col_reg}>=20'b00000110011001101001) && ({row_reg, col_reg}<20'b00000110100100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00000110100100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00000110100100011111) && ({row_reg, col_reg}<20'b00000110100101001000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00000110100101001000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00000110100101001001) && ({row_reg, col_reg}<20'b00000110100101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00000110100101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00000110100101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00000110100101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00000110100101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00000110100101010000) && ({row_reg, col_reg}<20'b00000110101000110111)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00000110101000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00000110101000111000) && ({row_reg, col_reg}<20'b00000110101000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00000110101000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00000110101000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00000110101000111100) && ({row_reg, col_reg}<20'b00000110101000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00000110101000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00000110101000111111) && ({row_reg, col_reg}<20'b00000110101001100001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00000110101001100001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00000110101001100010) && ({row_reg, col_reg}<20'b00000110101001100100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00000110101001100100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00000110101001100101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00000110101001100110) && ({row_reg, col_reg}<20'b00000110101001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00000110101001101000)) color_data = 12'b101110111011;

		if(({row_reg, col_reg}>=20'b00000110101001101001) && ({row_reg, col_reg}<20'b00000110110100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00000110110100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00000110110100011111) && ({row_reg, col_reg}<20'b00000110110101001000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00000110110101001000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00000110110101001001) && ({row_reg, col_reg}<20'b00000110110101001110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00000110110101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00000110110101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00000110110101010000) && ({row_reg, col_reg}<20'b00000110111000110111)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00000110111000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00000110111000111000) && ({row_reg, col_reg}<20'b00000110111000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00000110111000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00000110111000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00000110111000111100) && ({row_reg, col_reg}<20'b00000110111000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00000110111000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00000110111000111111) && ({row_reg, col_reg}<20'b00000110111001100001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00000110111001100001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00000110111001100010) && ({row_reg, col_reg}<20'b00000110111001100100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00000110111001100100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00000110111001100101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00000110111001100110) && ({row_reg, col_reg}<20'b00000110111001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00000110111001101000)) color_data = 12'b101110111011;

		if(({row_reg, col_reg}>=20'b00000110111001101001) && ({row_reg, col_reg}<20'b00000111000100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00000111000100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00000111000100011111) && ({row_reg, col_reg}<20'b00000111000101001110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00000111000101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00000111000101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00000111000101010000) && ({row_reg, col_reg}<20'b00000111001000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00000111001000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00000111001000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00000111001000111000) && ({row_reg, col_reg}<20'b00000111001000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00000111001000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00000111001000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00000111001000111100) && ({row_reg, col_reg}<20'b00000111001000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00000111001000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00000111001000111111) && ({row_reg, col_reg}<20'b00000111001001100001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00000111001001100001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00000111001001100010) && ({row_reg, col_reg}<20'b00000111001001100100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00000111001001100100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00000111001001100101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00000111001001100110) && ({row_reg, col_reg}<20'b00000111001001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00000111001001101000)) color_data = 12'b101110111011;

		if(({row_reg, col_reg}>=20'b00000111001001101001) && ({row_reg, col_reg}<20'b00000111010100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00000111010100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00000111010100011111) && ({row_reg, col_reg}<20'b00000111010101001110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00000111010101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00000111010101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00000111010101010000) && ({row_reg, col_reg}<20'b00000111011000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00000111011000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00000111011000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00000111011000111000) && ({row_reg, col_reg}<20'b00000111011000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00000111011000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00000111011000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00000111011000111100) && ({row_reg, col_reg}<20'b00000111011000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00000111011000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00000111011000111111) && ({row_reg, col_reg}<20'b00000111011001100001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00000111011001100001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00000111011001100010) && ({row_reg, col_reg}<20'b00000111011001100100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00000111011001100100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00000111011001100101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00000111011001100110) && ({row_reg, col_reg}<20'b00000111011001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00000111011001101000)) color_data = 12'b101110111011;

		if(({row_reg, col_reg}>=20'b00000111011001101001) && ({row_reg, col_reg}<20'b00000111100100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00000111100100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00000111100100011111) && ({row_reg, col_reg}<20'b00000111100101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00000111100101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00000111100101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00000111100101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00000111100101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00000111100101010000) && ({row_reg, col_reg}<20'b00000111101000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00000111101000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00000111101000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00000111101000111000) && ({row_reg, col_reg}<20'b00000111101000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00000111101000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00000111101000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00000111101000111100) && ({row_reg, col_reg}<20'b00000111101000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00000111101000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00000111101000111111) && ({row_reg, col_reg}<20'b00000111101001100001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00000111101001100001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00000111101001100010) && ({row_reg, col_reg}<20'b00000111101001100100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00000111101001100100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00000111101001100101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00000111101001100110) && ({row_reg, col_reg}<20'b00000111101001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00000111101001101000)) color_data = 12'b101110111011;

		if(({row_reg, col_reg}>=20'b00000111101001101001) && ({row_reg, col_reg}<20'b00000111110100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00000111110100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00000111110100011111) && ({row_reg, col_reg}<20'b00000111110101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00000111110101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00000111110101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00000111110101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00000111110101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00000111110101010000) && ({row_reg, col_reg}<20'b00000111111000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00000111111000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00000111111000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00000111111000111000) && ({row_reg, col_reg}<20'b00000111111000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00000111111000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00000111111000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00000111111000111100) && ({row_reg, col_reg}<20'b00000111111000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00000111111000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00000111111000111111) && ({row_reg, col_reg}<20'b00000111111001100100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00000111111001100100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00000111111001100101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00000111111001100110) && ({row_reg, col_reg}<20'b00000111111001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00000111111001101000)) color_data = 12'b101110111011;

		if(({row_reg, col_reg}>=20'b00000111111001101001) && ({row_reg, col_reg}<20'b00001000000100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00001000000100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00001000000100011111) && ({row_reg, col_reg}<20'b00001000000101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00001000000101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00001000000101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00001000000101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00001000000101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00001000000101010000) && ({row_reg, col_reg}<20'b00001000001000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00001000001000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00001000001000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00001000001000111000) && ({row_reg, col_reg}<20'b00001000001000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00001000001000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00001000001000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00001000001000111100) && ({row_reg, col_reg}<20'b00001000001000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00001000001000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00001000001000111111) && ({row_reg, col_reg}<20'b00001000001001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00001000001001100110) && ({row_reg, col_reg}<20'b00001000001001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00001000001001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00001000001001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00001000001001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00001000001001101011) && ({row_reg, col_reg}<20'b00001000010100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00001000010100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00001000010100011111) && ({row_reg, col_reg}<20'b00001000010101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00001000010101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00001000010101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00001000010101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00001000010101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00001000010101010000) && ({row_reg, col_reg}<20'b00001000011000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00001000011000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00001000011000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00001000011000111000) && ({row_reg, col_reg}<20'b00001000011000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00001000011000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00001000011000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00001000011000111100) && ({row_reg, col_reg}<20'b00001000011000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00001000011000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00001000011000111111) && ({row_reg, col_reg}<20'b00001000011001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00001000011001100110) && ({row_reg, col_reg}<20'b00001000011001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00001000011001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00001000011001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00001000011001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00001000011001101011) && ({row_reg, col_reg}<20'b00001000100100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00001000100100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00001000100100011111) && ({row_reg, col_reg}<20'b00001000100101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00001000100101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00001000100101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00001000100101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00001000100101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00001000100101010000) && ({row_reg, col_reg}<20'b00001000101000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00001000101000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00001000101000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00001000101000111000) && ({row_reg, col_reg}<20'b00001000101000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00001000101000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00001000101000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00001000101000111100) && ({row_reg, col_reg}<20'b00001000101000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00001000101000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00001000101000111111) && ({row_reg, col_reg}<20'b00001000101001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00001000101001100110) && ({row_reg, col_reg}<20'b00001000101001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00001000101001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00001000101001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00001000101001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00001000101001101011) && ({row_reg, col_reg}<20'b00001000110100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00001000110100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00001000110100011111) && ({row_reg, col_reg}<20'b00001000110101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00001000110101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00001000110101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00001000110101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00001000110101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00001000110101010000) && ({row_reg, col_reg}<20'b00001000111000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00001000111000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00001000111000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00001000111000111000) && ({row_reg, col_reg}<20'b00001000111000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00001000111000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00001000111000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00001000111000111100) && ({row_reg, col_reg}<20'b00001000111000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00001000111000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00001000111000111111) && ({row_reg, col_reg}<20'b00001000111001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00001000111001100110) && ({row_reg, col_reg}<20'b00001000111001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00001000111001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00001000111001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00001000111001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00001000111001101011) && ({row_reg, col_reg}<20'b00001001000100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00001001000100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00001001000100011111) && ({row_reg, col_reg}<20'b00001001000101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00001001000101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00001001000101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00001001000101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00001001000101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00001001000101010000) && ({row_reg, col_reg}<20'b00001001001000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00001001001000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00001001001000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00001001001000111000) && ({row_reg, col_reg}<20'b00001001001000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00001001001000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00001001001000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00001001001000111100) && ({row_reg, col_reg}<20'b00001001001000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00001001001000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00001001001000111111) && ({row_reg, col_reg}<20'b00001001001001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00001001001001100110) && ({row_reg, col_reg}<20'b00001001001001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00001001001001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00001001001001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00001001001001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00001001001001101011) && ({row_reg, col_reg}<20'b00001001010100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00001001010100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00001001010100011111) && ({row_reg, col_reg}<20'b00001001010101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00001001010101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00001001010101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00001001010101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00001001010101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00001001010101010000) && ({row_reg, col_reg}<20'b00001001011000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00001001011000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00001001011000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00001001011000111000) && ({row_reg, col_reg}<20'b00001001011000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00001001011000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00001001011000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00001001011000111100) && ({row_reg, col_reg}<20'b00001001011000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00001001011000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00001001011000111111) && ({row_reg, col_reg}<20'b00001001011001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00001001011001100110) && ({row_reg, col_reg}<20'b00001001011001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00001001011001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00001001011001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00001001011001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00001001011001101011) && ({row_reg, col_reg}<20'b00001001100100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00001001100100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00001001100100011111) && ({row_reg, col_reg}<20'b00001001100101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00001001100101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00001001100101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00001001100101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00001001100101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00001001100101010000) && ({row_reg, col_reg}<20'b00001001101000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00001001101000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00001001101000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00001001101000111000) && ({row_reg, col_reg}<20'b00001001101000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00001001101000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00001001101000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00001001101000111100) && ({row_reg, col_reg}<20'b00001001101000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00001001101000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00001001101000111111) && ({row_reg, col_reg}<20'b00001001101001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00001001101001100110) && ({row_reg, col_reg}<20'b00001001101001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00001001101001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00001001101001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00001001101001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00001001101001101011) && ({row_reg, col_reg}<20'b00001001110100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00001001110100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00001001110100011111) && ({row_reg, col_reg}<20'b00001001110101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00001001110101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00001001110101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00001001110101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00001001110101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00001001110101010000) && ({row_reg, col_reg}<20'b00001001111000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00001001111000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00001001111000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00001001111000111000) && ({row_reg, col_reg}<20'b00001001111000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00001001111000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00001001111000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00001001111000111100) && ({row_reg, col_reg}<20'b00001001111000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00001001111000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00001001111000111111) && ({row_reg, col_reg}<20'b00001001111001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00001001111001100110) && ({row_reg, col_reg}<20'b00001001111001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00001001111001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00001001111001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00001001111001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00001001111001101011) && ({row_reg, col_reg}<20'b00001010000100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00001010000100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00001010000100011111) && ({row_reg, col_reg}<20'b00001010000101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00001010000101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00001010000101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00001010000101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00001010000101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00001010000101010000) && ({row_reg, col_reg}<20'b00001010001000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00001010001000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00001010001000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00001010001000111000) && ({row_reg, col_reg}<20'b00001010001000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00001010001000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00001010001000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00001010001000111100) && ({row_reg, col_reg}<20'b00001010001000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00001010001000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00001010001000111111) && ({row_reg, col_reg}<20'b00001010001001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00001010001001100110) && ({row_reg, col_reg}<20'b00001010001001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00001010001001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00001010001001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00001010001001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00001010001001101011) && ({row_reg, col_reg}<20'b00001010010100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00001010010100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00001010010100011111) && ({row_reg, col_reg}<20'b00001010010101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00001010010101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00001010010101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00001010010101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00001010010101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00001010010101010000) && ({row_reg, col_reg}<20'b00001010011000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00001010011000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00001010011000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00001010011000111000) && ({row_reg, col_reg}<20'b00001010011000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00001010011000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00001010011000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00001010011000111100) && ({row_reg, col_reg}<20'b00001010011000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00001010011000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00001010011000111111) && ({row_reg, col_reg}<20'b00001010011001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00001010011001100110) && ({row_reg, col_reg}<20'b00001010011001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00001010011001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00001010011001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00001010011001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00001010011001101011) && ({row_reg, col_reg}<20'b00001010100100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00001010100100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00001010100100011111) && ({row_reg, col_reg}<20'b00001010100101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00001010100101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00001010100101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00001010100101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00001010100101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00001010100101010000) && ({row_reg, col_reg}<20'b00001010101000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00001010101000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00001010101000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00001010101000111000) && ({row_reg, col_reg}<20'b00001010101000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00001010101000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00001010101000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00001010101000111100) && ({row_reg, col_reg}<20'b00001010101000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00001010101000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00001010101000111111) && ({row_reg, col_reg}<20'b00001010101001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00001010101001100110) && ({row_reg, col_reg}<20'b00001010101001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00001010101001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00001010101001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00001010101001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00001010101001101011) && ({row_reg, col_reg}<20'b00001010110100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00001010110100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00001010110100011111) && ({row_reg, col_reg}<20'b00001010110101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00001010110101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00001010110101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00001010110101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00001010110101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00001010110101010000) && ({row_reg, col_reg}<20'b00001010111000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00001010111000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00001010111000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00001010111000111000) && ({row_reg, col_reg}<20'b00001010111000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00001010111000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00001010111000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00001010111000111100) && ({row_reg, col_reg}<20'b00001010111000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00001010111000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00001010111000111111) && ({row_reg, col_reg}<20'b00001010111001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00001010111001100110) && ({row_reg, col_reg}<20'b00001010111001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00001010111001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00001010111001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00001010111001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00001010111001101011) && ({row_reg, col_reg}<20'b00001011000100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00001011000100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00001011000100011111) && ({row_reg, col_reg}<20'b00001011000101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00001011000101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00001011000101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00001011000101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00001011000101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00001011000101010000) && ({row_reg, col_reg}<20'b00001011001000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00001011001000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00001011001000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00001011001000111000) && ({row_reg, col_reg}<20'b00001011001000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00001011001000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00001011001000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00001011001000111100) && ({row_reg, col_reg}<20'b00001011001000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00001011001000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00001011001000111111) && ({row_reg, col_reg}<20'b00001011001001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00001011001001100110) && ({row_reg, col_reg}<20'b00001011001001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00001011001001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00001011001001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00001011001001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00001011001001101011) && ({row_reg, col_reg}<20'b00001011010100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00001011010100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00001011010100011111) && ({row_reg, col_reg}<20'b00001011010101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00001011010101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00001011010101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00001011010101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00001011010101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00001011010101010000) && ({row_reg, col_reg}<20'b00001011011000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00001011011000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00001011011000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00001011011000111000) && ({row_reg, col_reg}<20'b00001011011000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00001011011000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00001011011000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00001011011000111100) && ({row_reg, col_reg}<20'b00001011011000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00001011011000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00001011011000111111) && ({row_reg, col_reg}<20'b00001011011001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00001011011001100110) && ({row_reg, col_reg}<20'b00001011011001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00001011011001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00001011011001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00001011011001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00001011011001101011) && ({row_reg, col_reg}<20'b00001011100100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00001011100100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00001011100100011111) && ({row_reg, col_reg}<20'b00001011100101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00001011100101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00001011100101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00001011100101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00001011100101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00001011100101010000) && ({row_reg, col_reg}<20'b00001011101000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00001011101000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00001011101000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00001011101000111000) && ({row_reg, col_reg}<20'b00001011101000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00001011101000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00001011101000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00001011101000111100) && ({row_reg, col_reg}<20'b00001011101000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00001011101000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00001011101000111111) && ({row_reg, col_reg}<20'b00001011101001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00001011101001100110) && ({row_reg, col_reg}<20'b00001011101001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00001011101001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00001011101001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00001011101001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00001011101001101011) && ({row_reg, col_reg}<20'b00001011110100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00001011110100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00001011110100011111) && ({row_reg, col_reg}<20'b00001011110101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00001011110101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00001011110101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00001011110101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00001011110101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00001011110101010000) && ({row_reg, col_reg}<20'b00001011111000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00001011111000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00001011111000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00001011111000111000) && ({row_reg, col_reg}<20'b00001011111000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00001011111000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00001011111000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00001011111000111100) && ({row_reg, col_reg}<20'b00001011111000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00001011111000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00001011111000111111) && ({row_reg, col_reg}<20'b00001011111001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00001011111001100110) && ({row_reg, col_reg}<20'b00001011111001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00001011111001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00001011111001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00001011111001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00001011111001101011) && ({row_reg, col_reg}<20'b00001100000100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00001100000100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00001100000100011111) && ({row_reg, col_reg}<20'b00001100000101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00001100000101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00001100000101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00001100000101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00001100000101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00001100000101010000) && ({row_reg, col_reg}<20'b00001100001000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00001100001000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00001100001000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00001100001000111000) && ({row_reg, col_reg}<20'b00001100001000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00001100001000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00001100001000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00001100001000111100) && ({row_reg, col_reg}<20'b00001100001000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00001100001000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00001100001000111111) && ({row_reg, col_reg}<20'b00001100001001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00001100001001100110) && ({row_reg, col_reg}<20'b00001100001001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00001100001001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00001100001001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00001100001001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00001100001001101011) && ({row_reg, col_reg}<20'b00001100010100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00001100010100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00001100010100011111) && ({row_reg, col_reg}<20'b00001100010101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00001100010101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00001100010101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00001100010101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00001100010101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00001100010101010000) && ({row_reg, col_reg}<20'b00001100011000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00001100011000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00001100011000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00001100011000111000) && ({row_reg, col_reg}<20'b00001100011000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00001100011000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00001100011000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00001100011000111100) && ({row_reg, col_reg}<20'b00001100011000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00001100011000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00001100011000111111) && ({row_reg, col_reg}<20'b00001100011001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00001100011001100110) && ({row_reg, col_reg}<20'b00001100011001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00001100011001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00001100011001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00001100011001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00001100011001101011) && ({row_reg, col_reg}<20'b00001100100100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00001100100100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00001100100100011111) && ({row_reg, col_reg}<20'b00001100100101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00001100100101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00001100100101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00001100100101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00001100100101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00001100100101010000) && ({row_reg, col_reg}<20'b00001100101000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00001100101000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00001100101000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00001100101000111000) && ({row_reg, col_reg}<20'b00001100101000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00001100101000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00001100101000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00001100101000111100) && ({row_reg, col_reg}<20'b00001100101000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00001100101000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00001100101000111111) && ({row_reg, col_reg}<20'b00001100101001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00001100101001100110) && ({row_reg, col_reg}<20'b00001100101001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00001100101001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00001100101001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00001100101001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00001100101001101011) && ({row_reg, col_reg}<20'b00001100110100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00001100110100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00001100110100011111) && ({row_reg, col_reg}<20'b00001100110101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00001100110101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00001100110101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00001100110101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00001100110101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00001100110101010000) && ({row_reg, col_reg}<20'b00001100111000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00001100111000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00001100111000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00001100111000111000) && ({row_reg, col_reg}<20'b00001100111000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00001100111000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00001100111000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00001100111000111100) && ({row_reg, col_reg}<20'b00001100111000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00001100111000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00001100111000111111) && ({row_reg, col_reg}<20'b00001100111001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00001100111001100110) && ({row_reg, col_reg}<20'b00001100111001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00001100111001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00001100111001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00001100111001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00001100111001101011) && ({row_reg, col_reg}<20'b00001101000100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00001101000100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00001101000100011111) && ({row_reg, col_reg}<20'b00001101000101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00001101000101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00001101000101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00001101000101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00001101000101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00001101000101010000) && ({row_reg, col_reg}<20'b00001101001000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00001101001000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00001101001000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00001101001000111000) && ({row_reg, col_reg}<20'b00001101001000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00001101001000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00001101001000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00001101001000111100) && ({row_reg, col_reg}<20'b00001101001000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00001101001000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00001101001000111111) && ({row_reg, col_reg}<20'b00001101001001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00001101001001100110) && ({row_reg, col_reg}<20'b00001101001001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00001101001001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00001101001001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00001101001001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00001101001001101011) && ({row_reg, col_reg}<20'b00001101010100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00001101010100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00001101010100011111) && ({row_reg, col_reg}<20'b00001101010101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00001101010101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00001101010101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00001101010101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00001101010101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00001101010101010000) && ({row_reg, col_reg}<20'b00001101011000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00001101011000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00001101011000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00001101011000111000) && ({row_reg, col_reg}<20'b00001101011000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00001101011000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00001101011000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00001101011000111100) && ({row_reg, col_reg}<20'b00001101011000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00001101011000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00001101011000111111) && ({row_reg, col_reg}<20'b00001101011001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00001101011001100110) && ({row_reg, col_reg}<20'b00001101011001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00001101011001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00001101011001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00001101011001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00001101011001101011) && ({row_reg, col_reg}<20'b00001101100100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00001101100100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00001101100100011111) && ({row_reg, col_reg}<20'b00001101100101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00001101100101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00001101100101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00001101100101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00001101100101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00001101100101010000) && ({row_reg, col_reg}<20'b00001101101000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00001101101000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00001101101000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00001101101000111000) && ({row_reg, col_reg}<20'b00001101101000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00001101101000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00001101101000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00001101101000111100) && ({row_reg, col_reg}<20'b00001101101000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00001101101000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00001101101000111111) && ({row_reg, col_reg}<20'b00001101101001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00001101101001100110) && ({row_reg, col_reg}<20'b00001101101001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00001101101001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00001101101001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00001101101001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00001101101001101011) && ({row_reg, col_reg}<20'b00001101110100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00001101110100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00001101110100011111) && ({row_reg, col_reg}<20'b00001101110101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00001101110101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00001101110101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00001101110101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00001101110101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00001101110101010000) && ({row_reg, col_reg}<20'b00001101111000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00001101111000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00001101111000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00001101111000111000) && ({row_reg, col_reg}<20'b00001101111000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00001101111000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00001101111000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00001101111000111100) && ({row_reg, col_reg}<20'b00001101111000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00001101111000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00001101111000111111) && ({row_reg, col_reg}<20'b00001101111001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00001101111001100110) && ({row_reg, col_reg}<20'b00001101111001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00001101111001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00001101111001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00001101111001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00001101111001101011) && ({row_reg, col_reg}<20'b00001110000100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00001110000100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00001110000100011111) && ({row_reg, col_reg}<20'b00001110000101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00001110000101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00001110000101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00001110000101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00001110000101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00001110000101010000) && ({row_reg, col_reg}<20'b00001110001000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00001110001000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00001110001000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00001110001000111000) && ({row_reg, col_reg}<20'b00001110001000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00001110001000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00001110001000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00001110001000111100) && ({row_reg, col_reg}<20'b00001110001000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00001110001000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00001110001000111111) && ({row_reg, col_reg}<20'b00001110001001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00001110001001100110) && ({row_reg, col_reg}<20'b00001110001001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00001110001001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00001110001001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00001110001001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00001110001001101011) && ({row_reg, col_reg}<20'b00001110010100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00001110010100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00001110010100011111) && ({row_reg, col_reg}<20'b00001110010101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00001110010101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00001110010101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00001110010101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00001110010101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00001110010101010000) && ({row_reg, col_reg}<20'b00001110011000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00001110011000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00001110011000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00001110011000111000) && ({row_reg, col_reg}<20'b00001110011000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00001110011000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00001110011000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00001110011000111100) && ({row_reg, col_reg}<20'b00001110011000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00001110011000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00001110011000111111) && ({row_reg, col_reg}<20'b00001110011001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00001110011001100110) && ({row_reg, col_reg}<20'b00001110011001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00001110011001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00001110011001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00001110011001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00001110011001101011) && ({row_reg, col_reg}<20'b00001110100100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00001110100100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00001110100100011111) && ({row_reg, col_reg}<20'b00001110100101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00001110100101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00001110100101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00001110100101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00001110100101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00001110100101010000) && ({row_reg, col_reg}<20'b00001110101000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00001110101000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00001110101000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00001110101000111000) && ({row_reg, col_reg}<20'b00001110101000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00001110101000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00001110101000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00001110101000111100) && ({row_reg, col_reg}<20'b00001110101000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00001110101000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00001110101000111111) && ({row_reg, col_reg}<20'b00001110101001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00001110101001100110) && ({row_reg, col_reg}<20'b00001110101001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00001110101001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00001110101001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00001110101001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00001110101001101011) && ({row_reg, col_reg}<20'b00001110110100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00001110110100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00001110110100011111) && ({row_reg, col_reg}<20'b00001110110101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00001110110101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00001110110101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00001110110101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00001110110101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00001110110101010000) && ({row_reg, col_reg}<20'b00001110111000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00001110111000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00001110111000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00001110111000111000) && ({row_reg, col_reg}<20'b00001110111000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00001110111000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00001110111000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00001110111000111100) && ({row_reg, col_reg}<20'b00001110111000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00001110111000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00001110111000111111) && ({row_reg, col_reg}<20'b00001110111001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00001110111001100110) && ({row_reg, col_reg}<20'b00001110111001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00001110111001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00001110111001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00001110111001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00001110111001101011) && ({row_reg, col_reg}<20'b00001111000100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00001111000100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00001111000100011111) && ({row_reg, col_reg}<20'b00001111000101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00001111000101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00001111000101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00001111000101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00001111000101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00001111000101010000) && ({row_reg, col_reg}<20'b00001111001000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00001111001000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00001111001000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00001111001000111000) && ({row_reg, col_reg}<20'b00001111001000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00001111001000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00001111001000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00001111001000111100) && ({row_reg, col_reg}<20'b00001111001000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00001111001000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00001111001000111111) && ({row_reg, col_reg}<20'b00001111001001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00001111001001100110) && ({row_reg, col_reg}<20'b00001111001001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00001111001001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00001111001001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00001111001001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00001111001001101011) && ({row_reg, col_reg}<20'b00001111010100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00001111010100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00001111010100011111) && ({row_reg, col_reg}<20'b00001111010101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00001111010101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00001111010101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00001111010101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00001111010101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00001111010101010000) && ({row_reg, col_reg}<20'b00001111011000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00001111011000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00001111011000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00001111011000111000) && ({row_reg, col_reg}<20'b00001111011000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00001111011000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00001111011000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00001111011000111100) && ({row_reg, col_reg}<20'b00001111011000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00001111011000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00001111011000111111) && ({row_reg, col_reg}<20'b00001111011001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00001111011001100110) && ({row_reg, col_reg}<20'b00001111011001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00001111011001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00001111011001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00001111011001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00001111011001101011) && ({row_reg, col_reg}<20'b00001111100100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00001111100100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00001111100100011111) && ({row_reg, col_reg}<20'b00001111100101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00001111100101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00001111100101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00001111100101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00001111100101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00001111100101010000) && ({row_reg, col_reg}<20'b00001111101000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00001111101000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00001111101000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00001111101000111000) && ({row_reg, col_reg}<20'b00001111101000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00001111101000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00001111101000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00001111101000111100) && ({row_reg, col_reg}<20'b00001111101000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00001111101000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00001111101000111111) && ({row_reg, col_reg}<20'b00001111101001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00001111101001100110) && ({row_reg, col_reg}<20'b00001111101001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00001111101001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00001111101001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00001111101001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00001111101001101011) && ({row_reg, col_reg}<20'b00001111110100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00001111110100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00001111110100011111) && ({row_reg, col_reg}<20'b00001111110101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00001111110101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00001111110101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00001111110101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00001111110101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00001111110101010000) && ({row_reg, col_reg}<20'b00001111111000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00001111111000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00001111111000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00001111111000111000) && ({row_reg, col_reg}<20'b00001111111000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00001111111000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00001111111000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00001111111000111100) && ({row_reg, col_reg}<20'b00001111111000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00001111111000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00001111111000111111) && ({row_reg, col_reg}<20'b00001111111001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00001111111001100110) && ({row_reg, col_reg}<20'b00001111111001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00001111111001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00001111111001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00001111111001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00001111111001101011) && ({row_reg, col_reg}<20'b00010000000100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00010000000100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00010000000100011111) && ({row_reg, col_reg}<20'b00010000000101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00010000000101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00010000000101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00010000000101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00010000000101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00010000000101010000) && ({row_reg, col_reg}<20'b00010000001000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00010000001000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00010000001000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00010000001000111000) && ({row_reg, col_reg}<20'b00010000001000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00010000001000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00010000001000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00010000001000111100) && ({row_reg, col_reg}<20'b00010000001000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00010000001000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00010000001000111111) && ({row_reg, col_reg}<20'b00010000001001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00010000001001100110) && ({row_reg, col_reg}<20'b00010000001001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00010000001001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00010000001001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00010000001001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00010000001001101011) && ({row_reg, col_reg}<20'b00010000010100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00010000010100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00010000010100011111) && ({row_reg, col_reg}<20'b00010000010101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00010000010101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00010000010101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00010000010101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00010000010101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00010000010101010000) && ({row_reg, col_reg}<20'b00010000011000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00010000011000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00010000011000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00010000011000111000) && ({row_reg, col_reg}<20'b00010000011000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00010000011000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00010000011000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00010000011000111100) && ({row_reg, col_reg}<20'b00010000011000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00010000011000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00010000011000111111) && ({row_reg, col_reg}<20'b00010000011001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00010000011001100110) && ({row_reg, col_reg}<20'b00010000011001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00010000011001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00010000011001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00010000011001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00010000011001101011) && ({row_reg, col_reg}<20'b00010000100100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00010000100100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00010000100100011111) && ({row_reg, col_reg}<20'b00010000100101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00010000100101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00010000100101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00010000100101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00010000100101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00010000100101010000) && ({row_reg, col_reg}<20'b00010000101000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00010000101000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00010000101000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00010000101000111000) && ({row_reg, col_reg}<20'b00010000101000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00010000101000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00010000101000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00010000101000111100) && ({row_reg, col_reg}<20'b00010000101000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00010000101000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00010000101000111111) && ({row_reg, col_reg}<20'b00010000101001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00010000101001100110) && ({row_reg, col_reg}<20'b00010000101001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00010000101001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00010000101001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00010000101001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00010000101001101011) && ({row_reg, col_reg}<20'b00010000110100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00010000110100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00010000110100011111) && ({row_reg, col_reg}<20'b00010000110101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00010000110101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00010000110101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00010000110101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00010000110101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00010000110101010000) && ({row_reg, col_reg}<20'b00010000111000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00010000111000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00010000111000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00010000111000111000) && ({row_reg, col_reg}<20'b00010000111000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00010000111000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00010000111000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00010000111000111100) && ({row_reg, col_reg}<20'b00010000111000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00010000111000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00010000111000111111) && ({row_reg, col_reg}<20'b00010000111001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00010000111001100110) && ({row_reg, col_reg}<20'b00010000111001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00010000111001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00010000111001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00010000111001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00010000111001101011) && ({row_reg, col_reg}<20'b00010001000100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00010001000100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00010001000100011111) && ({row_reg, col_reg}<20'b00010001000101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00010001000101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00010001000101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00010001000101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00010001000101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00010001000101010000) && ({row_reg, col_reg}<20'b00010001001000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00010001001000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00010001001000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00010001001000111000) && ({row_reg, col_reg}<20'b00010001001000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00010001001000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00010001001000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00010001001000111100) && ({row_reg, col_reg}<20'b00010001001000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00010001001000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00010001001000111111) && ({row_reg, col_reg}<20'b00010001001001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00010001001001100110) && ({row_reg, col_reg}<20'b00010001001001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00010001001001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00010001001001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00010001001001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00010001001001101011) && ({row_reg, col_reg}<20'b00010001010100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00010001010100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00010001010100011111) && ({row_reg, col_reg}<20'b00010001010101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00010001010101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00010001010101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00010001010101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00010001010101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00010001010101010000) && ({row_reg, col_reg}<20'b00010001011000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00010001011000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00010001011000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00010001011000111000) && ({row_reg, col_reg}<20'b00010001011000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00010001011000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00010001011000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00010001011000111100) && ({row_reg, col_reg}<20'b00010001011000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00010001011000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00010001011000111111) && ({row_reg, col_reg}<20'b00010001011001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00010001011001100110) && ({row_reg, col_reg}<20'b00010001011001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00010001011001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00010001011001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00010001011001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00010001011001101011) && ({row_reg, col_reg}<20'b00010001100100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00010001100100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00010001100100011111) && ({row_reg, col_reg}<20'b00010001100101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00010001100101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00010001100101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00010001100101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00010001100101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00010001100101010000) && ({row_reg, col_reg}<20'b00010001101000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00010001101000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00010001101000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00010001101000111000) && ({row_reg, col_reg}<20'b00010001101000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00010001101000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00010001101000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00010001101000111100) && ({row_reg, col_reg}<20'b00010001101000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00010001101000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00010001101000111111) && ({row_reg, col_reg}<20'b00010001101001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00010001101001100110) && ({row_reg, col_reg}<20'b00010001101001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00010001101001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00010001101001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00010001101001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00010001101001101011) && ({row_reg, col_reg}<20'b00010001110100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00010001110100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00010001110100011111) && ({row_reg, col_reg}<20'b00010001110101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00010001110101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00010001110101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00010001110101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00010001110101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00010001110101010000) && ({row_reg, col_reg}<20'b00010001111000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00010001111000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00010001111000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00010001111000111000) && ({row_reg, col_reg}<20'b00010001111000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00010001111000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00010001111000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00010001111000111100) && ({row_reg, col_reg}<20'b00010001111000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00010001111000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00010001111000111111) && ({row_reg, col_reg}<20'b00010001111001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00010001111001100110) && ({row_reg, col_reg}<20'b00010001111001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00010001111001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00010001111001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00010001111001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00010001111001101011) && ({row_reg, col_reg}<20'b00010010000100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00010010000100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00010010000100011111) && ({row_reg, col_reg}<20'b00010010000101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00010010000101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00010010000101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00010010000101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00010010000101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00010010000101010000) && ({row_reg, col_reg}<20'b00010010001000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00010010001000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00010010001000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00010010001000111000) && ({row_reg, col_reg}<20'b00010010001000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00010010001000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00010010001000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00010010001000111100) && ({row_reg, col_reg}<20'b00010010001000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00010010001000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00010010001000111111) && ({row_reg, col_reg}<20'b00010010001001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00010010001001100110) && ({row_reg, col_reg}<20'b00010010001001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00010010001001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00010010001001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00010010001001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00010010001001101011) && ({row_reg, col_reg}<20'b00010010010100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00010010010100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00010010010100011111) && ({row_reg, col_reg}<20'b00010010010101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00010010010101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00010010010101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00010010010101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00010010010101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00010010010101010000) && ({row_reg, col_reg}<20'b00010010011000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00010010011000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00010010011000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00010010011000111000) && ({row_reg, col_reg}<20'b00010010011000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00010010011000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00010010011000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00010010011000111100) && ({row_reg, col_reg}<20'b00010010011000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00010010011000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00010010011000111111) && ({row_reg, col_reg}<20'b00010010011001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00010010011001100110) && ({row_reg, col_reg}<20'b00010010011001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00010010011001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00010010011001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00010010011001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00010010011001101011) && ({row_reg, col_reg}<20'b00010010100100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00010010100100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00010010100100011111) && ({row_reg, col_reg}<20'b00010010100101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00010010100101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00010010100101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00010010100101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00010010100101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00010010100101010000) && ({row_reg, col_reg}<20'b00010010101000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00010010101000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00010010101000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00010010101000111000) && ({row_reg, col_reg}<20'b00010010101000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00010010101000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00010010101000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00010010101000111100) && ({row_reg, col_reg}<20'b00010010101000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00010010101000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00010010101000111111) && ({row_reg, col_reg}<20'b00010010101001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00010010101001100110) && ({row_reg, col_reg}<20'b00010010101001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00010010101001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00010010101001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00010010101001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00010010101001101011) && ({row_reg, col_reg}<20'b00010010110100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00010010110100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00010010110100011111) && ({row_reg, col_reg}<20'b00010010110101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00010010110101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00010010110101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00010010110101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00010010110101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00010010110101010000) && ({row_reg, col_reg}<20'b00010010111000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00010010111000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00010010111000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00010010111000111000) && ({row_reg, col_reg}<20'b00010010111000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00010010111000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00010010111000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00010010111000111100) && ({row_reg, col_reg}<20'b00010010111000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00010010111000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00010010111000111111) && ({row_reg, col_reg}<20'b00010010111001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00010010111001100110) && ({row_reg, col_reg}<20'b00010010111001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00010010111001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00010010111001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00010010111001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00010010111001101011) && ({row_reg, col_reg}<20'b00010011000100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00010011000100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00010011000100011111) && ({row_reg, col_reg}<20'b00010011000101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00010011000101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00010011000101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00010011000101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00010011000101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00010011000101010000) && ({row_reg, col_reg}<20'b00010011001000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00010011001000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00010011001000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00010011001000111000) && ({row_reg, col_reg}<20'b00010011001000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00010011001000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00010011001000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00010011001000111100) && ({row_reg, col_reg}<20'b00010011001000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00010011001000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00010011001000111111) && ({row_reg, col_reg}<20'b00010011001001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00010011001001100110) && ({row_reg, col_reg}<20'b00010011001001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00010011001001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00010011001001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00010011001001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00010011001001101011) && ({row_reg, col_reg}<20'b00010011010100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00010011010100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00010011010100011111) && ({row_reg, col_reg}<20'b00010011010101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00010011010101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00010011010101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00010011010101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00010011010101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00010011010101010000) && ({row_reg, col_reg}<20'b00010011011000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00010011011000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00010011011000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00010011011000111000) && ({row_reg, col_reg}<20'b00010011011000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00010011011000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00010011011000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00010011011000111100) && ({row_reg, col_reg}<20'b00010011011000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00010011011000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00010011011000111111) && ({row_reg, col_reg}<20'b00010011011001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00010011011001100110) && ({row_reg, col_reg}<20'b00010011011001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00010011011001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00010011011001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00010011011001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00010011011001101011) && ({row_reg, col_reg}<20'b00010011100100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00010011100100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00010011100100011111) && ({row_reg, col_reg}<20'b00010011100101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00010011100101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00010011100101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00010011100101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00010011100101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00010011100101010000) && ({row_reg, col_reg}<20'b00010011101000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00010011101000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00010011101000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00010011101000111000) && ({row_reg, col_reg}<20'b00010011101000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00010011101000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00010011101000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00010011101000111100) && ({row_reg, col_reg}<20'b00010011101000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00010011101000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00010011101000111111) && ({row_reg, col_reg}<20'b00010011101001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00010011101001100110) && ({row_reg, col_reg}<20'b00010011101001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00010011101001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00010011101001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00010011101001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00010011101001101011) && ({row_reg, col_reg}<20'b00010011110100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00010011110100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00010011110100011111) && ({row_reg, col_reg}<20'b00010011110101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00010011110101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00010011110101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00010011110101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00010011110101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00010011110101010000) && ({row_reg, col_reg}<20'b00010011111000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00010011111000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00010011111000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00010011111000111000) && ({row_reg, col_reg}<20'b00010011111000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00010011111000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00010011111000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00010011111000111100) && ({row_reg, col_reg}<20'b00010011111000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00010011111000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00010011111000111111) && ({row_reg, col_reg}<20'b00010011111001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00010011111001100110) && ({row_reg, col_reg}<20'b00010011111001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00010011111001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00010011111001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00010011111001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00010011111001101011) && ({row_reg, col_reg}<20'b00010100000100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00010100000100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00010100000100011111) && ({row_reg, col_reg}<20'b00010100000101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00010100000101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00010100000101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00010100000101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00010100000101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00010100000101010000) && ({row_reg, col_reg}<20'b00010100001000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00010100001000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00010100001000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00010100001000111000) && ({row_reg, col_reg}<20'b00010100001000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00010100001000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00010100001000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00010100001000111100) && ({row_reg, col_reg}<20'b00010100001000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00010100001000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00010100001000111111) && ({row_reg, col_reg}<20'b00010100001001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00010100001001100110) && ({row_reg, col_reg}<20'b00010100001001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00010100001001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00010100001001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00010100001001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00010100001001101011) && ({row_reg, col_reg}<20'b00010100010100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00010100010100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00010100010100011111) && ({row_reg, col_reg}<20'b00010100010101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00010100010101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00010100010101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00010100010101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00010100010101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00010100010101010000) && ({row_reg, col_reg}<20'b00010100011000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00010100011000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00010100011000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00010100011000111000) && ({row_reg, col_reg}<20'b00010100011000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00010100011000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00010100011000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00010100011000111100) && ({row_reg, col_reg}<20'b00010100011000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00010100011000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00010100011000111111) && ({row_reg, col_reg}<20'b00010100011001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00010100011001100110) && ({row_reg, col_reg}<20'b00010100011001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00010100011001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00010100011001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00010100011001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00010100011001101011) && ({row_reg, col_reg}<20'b00010100100100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00010100100100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00010100100100011111) && ({row_reg, col_reg}<20'b00010100100101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00010100100101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00010100100101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00010100100101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00010100100101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00010100100101010000) && ({row_reg, col_reg}<20'b00010100101000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00010100101000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00010100101000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00010100101000111000) && ({row_reg, col_reg}<20'b00010100101000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00010100101000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00010100101000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00010100101000111100) && ({row_reg, col_reg}<20'b00010100101000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00010100101000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00010100101000111111) && ({row_reg, col_reg}<20'b00010100101001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00010100101001100110) && ({row_reg, col_reg}<20'b00010100101001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00010100101001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00010100101001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00010100101001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00010100101001101011) && ({row_reg, col_reg}<20'b00010100110100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00010100110100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00010100110100011111) && ({row_reg, col_reg}<20'b00010100110101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00010100110101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00010100110101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00010100110101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00010100110101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00010100110101010000) && ({row_reg, col_reg}<20'b00010100111000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00010100111000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00010100111000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00010100111000111000) && ({row_reg, col_reg}<20'b00010100111000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00010100111000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00010100111000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00010100111000111100) && ({row_reg, col_reg}<20'b00010100111000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00010100111000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00010100111000111111) && ({row_reg, col_reg}<20'b00010100111001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00010100111001100110) && ({row_reg, col_reg}<20'b00010100111001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00010100111001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00010100111001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00010100111001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00010100111001101011) && ({row_reg, col_reg}<20'b00010101000100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00010101000100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00010101000100011111) && ({row_reg, col_reg}<20'b00010101000101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00010101000101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00010101000101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00010101000101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00010101000101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00010101000101010000) && ({row_reg, col_reg}<20'b00010101001000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00010101001000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00010101001000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00010101001000111000) && ({row_reg, col_reg}<20'b00010101001000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00010101001000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00010101001000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00010101001000111100) && ({row_reg, col_reg}<20'b00010101001000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00010101001000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00010101001000111111) && ({row_reg, col_reg}<20'b00010101001001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00010101001001100110) && ({row_reg, col_reg}<20'b00010101001001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00010101001001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00010101001001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00010101001001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00010101001001101011) && ({row_reg, col_reg}<20'b00010101010100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00010101010100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00010101010100011111) && ({row_reg, col_reg}<20'b00010101010101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00010101010101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00010101010101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00010101010101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00010101010101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00010101010101010000) && ({row_reg, col_reg}<20'b00010101011000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00010101011000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00010101011000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00010101011000111000) && ({row_reg, col_reg}<20'b00010101011000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00010101011000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00010101011000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00010101011000111100) && ({row_reg, col_reg}<20'b00010101011000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00010101011000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00010101011000111111) && ({row_reg, col_reg}<20'b00010101011001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00010101011001100110) && ({row_reg, col_reg}<20'b00010101011001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00010101011001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00010101011001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00010101011001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00010101011001101011) && ({row_reg, col_reg}<20'b00010101100100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00010101100100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00010101100100011111) && ({row_reg, col_reg}<20'b00010101100101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00010101100101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00010101100101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00010101100101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00010101100101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00010101100101010000) && ({row_reg, col_reg}<20'b00010101101000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00010101101000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00010101101000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00010101101000111000) && ({row_reg, col_reg}<20'b00010101101000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00010101101000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00010101101000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00010101101000111100) && ({row_reg, col_reg}<20'b00010101101000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00010101101000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00010101101000111111) && ({row_reg, col_reg}<20'b00010101101001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00010101101001100110) && ({row_reg, col_reg}<20'b00010101101001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00010101101001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00010101101001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00010101101001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00010101101001101011) && ({row_reg, col_reg}<20'b00010101110100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00010101110100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00010101110100011111) && ({row_reg, col_reg}<20'b00010101110101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00010101110101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00010101110101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00010101110101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00010101110101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00010101110101010000) && ({row_reg, col_reg}<20'b00010101111000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00010101111000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00010101111000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00010101111000111000) && ({row_reg, col_reg}<20'b00010101111000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00010101111000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00010101111000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00010101111000111100) && ({row_reg, col_reg}<20'b00010101111000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00010101111000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00010101111000111111) && ({row_reg, col_reg}<20'b00010101111001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00010101111001100110) && ({row_reg, col_reg}<20'b00010101111001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00010101111001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00010101111001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00010101111001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00010101111001101011) && ({row_reg, col_reg}<20'b00010110000100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00010110000100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00010110000100011111) && ({row_reg, col_reg}<20'b00010110000101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00010110000101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00010110000101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00010110000101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00010110000101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00010110000101010000) && ({row_reg, col_reg}<20'b00010110001000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00010110001000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00010110001000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00010110001000111000) && ({row_reg, col_reg}<20'b00010110001000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00010110001000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00010110001000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00010110001000111100) && ({row_reg, col_reg}<20'b00010110001000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00010110001000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00010110001000111111) && ({row_reg, col_reg}<20'b00010110001001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00010110001001100110) && ({row_reg, col_reg}<20'b00010110001001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00010110001001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00010110001001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00010110001001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00010110001001101011) && ({row_reg, col_reg}<20'b00010110010100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00010110010100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00010110010100011111) && ({row_reg, col_reg}<20'b00010110010101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00010110010101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00010110010101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00010110010101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00010110010101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00010110010101010000) && ({row_reg, col_reg}<20'b00010110011000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00010110011000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00010110011000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00010110011000111000) && ({row_reg, col_reg}<20'b00010110011000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00010110011000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00010110011000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00010110011000111100) && ({row_reg, col_reg}<20'b00010110011000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00010110011000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00010110011000111111) && ({row_reg, col_reg}<20'b00010110011001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00010110011001100110) && ({row_reg, col_reg}<20'b00010110011001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00010110011001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00010110011001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00010110011001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00010110011001101011) && ({row_reg, col_reg}<20'b00010110100100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00010110100100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00010110100100011111) && ({row_reg, col_reg}<20'b00010110100101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00010110100101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00010110100101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00010110100101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00010110100101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00010110100101010000) && ({row_reg, col_reg}<20'b00010110101000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00010110101000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00010110101000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00010110101000111000) && ({row_reg, col_reg}<20'b00010110101000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00010110101000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00010110101000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00010110101000111100) && ({row_reg, col_reg}<20'b00010110101000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00010110101000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00010110101000111111) && ({row_reg, col_reg}<20'b00010110101001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00010110101001100110) && ({row_reg, col_reg}<20'b00010110101001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00010110101001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00010110101001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00010110101001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00010110101001101011) && ({row_reg, col_reg}<20'b00010110110100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00010110110100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00010110110100011111) && ({row_reg, col_reg}<20'b00010110110101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00010110110101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00010110110101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00010110110101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00010110110101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00010110110101010000) && ({row_reg, col_reg}<20'b00010110111000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00010110111000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00010110111000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00010110111000111000) && ({row_reg, col_reg}<20'b00010110111000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00010110111000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00010110111000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00010110111000111100) && ({row_reg, col_reg}<20'b00010110111000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00010110111000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00010110111000111111) && ({row_reg, col_reg}<20'b00010110111001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00010110111001100110) && ({row_reg, col_reg}<20'b00010110111001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00010110111001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00010110111001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00010110111001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00010110111001101011) && ({row_reg, col_reg}<20'b00010111000100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00010111000100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00010111000100011111) && ({row_reg, col_reg}<20'b00010111000101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00010111000101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00010111000101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00010111000101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00010111000101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00010111000101010000) && ({row_reg, col_reg}<20'b00010111001000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00010111001000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00010111001000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00010111001000111000) && ({row_reg, col_reg}<20'b00010111001000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00010111001000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00010111001000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00010111001000111100) && ({row_reg, col_reg}<20'b00010111001000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00010111001000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00010111001000111111) && ({row_reg, col_reg}<20'b00010111001001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00010111001001100110) && ({row_reg, col_reg}<20'b00010111001001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00010111001001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00010111001001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00010111001001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00010111001001101011) && ({row_reg, col_reg}<20'b00010111010100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00010111010100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00010111010100011111) && ({row_reg, col_reg}<20'b00010111010101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00010111010101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00010111010101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00010111010101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00010111010101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00010111010101010000) && ({row_reg, col_reg}<20'b00010111011000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00010111011000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00010111011000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00010111011000111000) && ({row_reg, col_reg}<20'b00010111011000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00010111011000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00010111011000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00010111011000111100) && ({row_reg, col_reg}<20'b00010111011000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00010111011000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00010111011000111111) && ({row_reg, col_reg}<20'b00010111011001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00010111011001100110) && ({row_reg, col_reg}<20'b00010111011001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00010111011001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00010111011001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00010111011001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00010111011001101011) && ({row_reg, col_reg}<20'b00010111100100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00010111100100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00010111100100011111) && ({row_reg, col_reg}<20'b00010111100101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00010111100101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00010111100101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00010111100101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00010111100101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00010111100101010000) && ({row_reg, col_reg}<20'b00010111101000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00010111101000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00010111101000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00010111101000111000) && ({row_reg, col_reg}<20'b00010111101000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00010111101000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00010111101000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00010111101000111100) && ({row_reg, col_reg}<20'b00010111101000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00010111101000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00010111101000111111) && ({row_reg, col_reg}<20'b00010111101001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00010111101001100110) && ({row_reg, col_reg}<20'b00010111101001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00010111101001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00010111101001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00010111101001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00010111101001101011) && ({row_reg, col_reg}<20'b00010111110100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00010111110100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00010111110100011111) && ({row_reg, col_reg}<20'b00010111110101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00010111110101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00010111110101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00010111110101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00010111110101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00010111110101010000) && ({row_reg, col_reg}<20'b00010111111000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00010111111000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00010111111000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00010111111000111000) && ({row_reg, col_reg}<20'b00010111111000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00010111111000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00010111111000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00010111111000111100) && ({row_reg, col_reg}<20'b00010111111000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00010111111000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00010111111000111111) && ({row_reg, col_reg}<20'b00010111111001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00010111111001100110) && ({row_reg, col_reg}<20'b00010111111001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00010111111001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00010111111001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00010111111001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00010111111001101011) && ({row_reg, col_reg}<20'b00011000000100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00011000000100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00011000000100011111) && ({row_reg, col_reg}<20'b00011000000101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00011000000101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00011000000101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00011000000101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00011000000101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00011000000101010000) && ({row_reg, col_reg}<20'b00011000001000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00011000001000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00011000001000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00011000001000111000) && ({row_reg, col_reg}<20'b00011000001000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00011000001000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00011000001000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00011000001000111100) && ({row_reg, col_reg}<20'b00011000001000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00011000001000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00011000001000111111) && ({row_reg, col_reg}<20'b00011000001001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00011000001001100110) && ({row_reg, col_reg}<20'b00011000001001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00011000001001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00011000001001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00011000001001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00011000001001101011) && ({row_reg, col_reg}<20'b00011000010100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00011000010100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00011000010100011111) && ({row_reg, col_reg}<20'b00011000010101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00011000010101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00011000010101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00011000010101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00011000010101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00011000010101010000) && ({row_reg, col_reg}<20'b00011000011000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00011000011000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00011000011000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00011000011000111000) && ({row_reg, col_reg}<20'b00011000011000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00011000011000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00011000011000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00011000011000111100) && ({row_reg, col_reg}<20'b00011000011000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00011000011000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00011000011000111111) && ({row_reg, col_reg}<20'b00011000011001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00011000011001100110) && ({row_reg, col_reg}<20'b00011000011001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00011000011001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00011000011001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00011000011001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00011000011001101011) && ({row_reg, col_reg}<20'b00011000100100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00011000100100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00011000100100011111) && ({row_reg, col_reg}<20'b00011000100101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00011000100101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00011000100101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00011000100101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00011000100101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00011000100101010000) && ({row_reg, col_reg}<20'b00011000101000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00011000101000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00011000101000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00011000101000111000) && ({row_reg, col_reg}<20'b00011000101000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00011000101000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00011000101000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00011000101000111100) && ({row_reg, col_reg}<20'b00011000101000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00011000101000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00011000101000111111) && ({row_reg, col_reg}<20'b00011000101001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00011000101001100110) && ({row_reg, col_reg}<20'b00011000101001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00011000101001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00011000101001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00011000101001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00011000101001101011) && ({row_reg, col_reg}<20'b00011000110100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00011000110100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00011000110100011111) && ({row_reg, col_reg}<20'b00011000110101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00011000110101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00011000110101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00011000110101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00011000110101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00011000110101010000) && ({row_reg, col_reg}<20'b00011000111000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00011000111000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00011000111000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00011000111000111000) && ({row_reg, col_reg}<20'b00011000111000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00011000111000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00011000111000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00011000111000111100) && ({row_reg, col_reg}<20'b00011000111000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00011000111000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00011000111000111111) && ({row_reg, col_reg}<20'b00011000111001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00011000111001100110) && ({row_reg, col_reg}<20'b00011000111001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00011000111001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00011000111001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00011000111001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00011000111001101011) && ({row_reg, col_reg}<20'b00011001000100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00011001000100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00011001000100011111) && ({row_reg, col_reg}<20'b00011001000101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00011001000101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00011001000101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00011001000101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00011001000101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00011001000101010000) && ({row_reg, col_reg}<20'b00011001001000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00011001001000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00011001001000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00011001001000111000) && ({row_reg, col_reg}<20'b00011001001000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00011001001000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00011001001000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00011001001000111100) && ({row_reg, col_reg}<20'b00011001001000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00011001001000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00011001001000111111) && ({row_reg, col_reg}<20'b00011001001001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00011001001001100110) && ({row_reg, col_reg}<20'b00011001001001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00011001001001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00011001001001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00011001001001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00011001001001101011) && ({row_reg, col_reg}<20'b00011001010100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00011001010100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00011001010100011111) && ({row_reg, col_reg}<20'b00011001010101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00011001010101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00011001010101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00011001010101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00011001010101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00011001010101010000) && ({row_reg, col_reg}<20'b00011001011000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00011001011000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00011001011000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00011001011000111000) && ({row_reg, col_reg}<20'b00011001011000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00011001011000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00011001011000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00011001011000111100) && ({row_reg, col_reg}<20'b00011001011000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00011001011000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00011001011000111111) && ({row_reg, col_reg}<20'b00011001011001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00011001011001100110) && ({row_reg, col_reg}<20'b00011001011001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00011001011001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00011001011001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00011001011001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00011001011001101011) && ({row_reg, col_reg}<20'b00011001100100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00011001100100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00011001100100011111) && ({row_reg, col_reg}<20'b00011001100101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00011001100101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00011001100101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00011001100101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00011001100101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00011001100101010000) && ({row_reg, col_reg}<20'b00011001101000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00011001101000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00011001101000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00011001101000111000) && ({row_reg, col_reg}<20'b00011001101000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00011001101000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00011001101000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00011001101000111100) && ({row_reg, col_reg}<20'b00011001101000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00011001101000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00011001101000111111) && ({row_reg, col_reg}<20'b00011001101001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00011001101001100110) && ({row_reg, col_reg}<20'b00011001101001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00011001101001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00011001101001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00011001101001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00011001101001101011) && ({row_reg, col_reg}<20'b00011001110100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00011001110100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00011001110100011111) && ({row_reg, col_reg}<20'b00011001110101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00011001110101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00011001110101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00011001110101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00011001110101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00011001110101010000) && ({row_reg, col_reg}<20'b00011001111000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00011001111000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00011001111000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00011001111000111000) && ({row_reg, col_reg}<20'b00011001111000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00011001111000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00011001111000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00011001111000111100) && ({row_reg, col_reg}<20'b00011001111000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00011001111000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00011001111000111111) && ({row_reg, col_reg}<20'b00011001111001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00011001111001100110) && ({row_reg, col_reg}<20'b00011001111001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00011001111001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00011001111001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00011001111001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00011001111001101011) && ({row_reg, col_reg}<20'b00011010000100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00011010000100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00011010000100011111) && ({row_reg, col_reg}<20'b00011010000101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00011010000101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00011010000101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00011010000101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00011010000101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00011010000101010000) && ({row_reg, col_reg}<20'b00011010001000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00011010001000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00011010001000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00011010001000111000) && ({row_reg, col_reg}<20'b00011010001000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00011010001000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00011010001000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00011010001000111100) && ({row_reg, col_reg}<20'b00011010001000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00011010001000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00011010001000111111) && ({row_reg, col_reg}<20'b00011010001001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00011010001001100110) && ({row_reg, col_reg}<20'b00011010001001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00011010001001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00011010001001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00011010001001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00011010001001101011) && ({row_reg, col_reg}<20'b00011010010100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00011010010100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00011010010100011111) && ({row_reg, col_reg}<20'b00011010010101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00011010010101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00011010010101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00011010010101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00011010010101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00011010010101010000) && ({row_reg, col_reg}<20'b00011010011000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00011010011000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00011010011000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00011010011000111000) && ({row_reg, col_reg}<20'b00011010011000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00011010011000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00011010011000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00011010011000111100) && ({row_reg, col_reg}<20'b00011010011000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00011010011000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00011010011000111111) && ({row_reg, col_reg}<20'b00011010011001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00011010011001100110) && ({row_reg, col_reg}<20'b00011010011001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00011010011001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00011010011001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00011010011001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00011010011001101011) && ({row_reg, col_reg}<20'b00011010100100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00011010100100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00011010100100011111) && ({row_reg, col_reg}<20'b00011010100101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00011010100101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00011010100101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00011010100101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00011010100101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00011010100101010000) && ({row_reg, col_reg}<20'b00011010101000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00011010101000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00011010101000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00011010101000111000) && ({row_reg, col_reg}<20'b00011010101000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00011010101000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00011010101000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00011010101000111100) && ({row_reg, col_reg}<20'b00011010101000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00011010101000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00011010101000111111) && ({row_reg, col_reg}<20'b00011010101001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00011010101001100110) && ({row_reg, col_reg}<20'b00011010101001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00011010101001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00011010101001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00011010101001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00011010101001101011) && ({row_reg, col_reg}<20'b00011010110100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00011010110100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00011010110100011111) && ({row_reg, col_reg}<20'b00011010110101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00011010110101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00011010110101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00011010110101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00011010110101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00011010110101010000) && ({row_reg, col_reg}<20'b00011010111000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00011010111000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00011010111000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00011010111000111000) && ({row_reg, col_reg}<20'b00011010111000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00011010111000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00011010111000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00011010111000111100) && ({row_reg, col_reg}<20'b00011010111000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00011010111000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00011010111000111111) && ({row_reg, col_reg}<20'b00011010111001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00011010111001100110) && ({row_reg, col_reg}<20'b00011010111001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00011010111001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00011010111001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00011010111001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00011010111001101011) && ({row_reg, col_reg}<20'b00011011000100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00011011000100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00011011000100011111) && ({row_reg, col_reg}<20'b00011011000101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00011011000101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00011011000101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00011011000101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00011011000101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00011011000101010000) && ({row_reg, col_reg}<20'b00011011001000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00011011001000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00011011001000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00011011001000111000) && ({row_reg, col_reg}<20'b00011011001000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00011011001000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00011011001000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00011011001000111100) && ({row_reg, col_reg}<20'b00011011001000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00011011001000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00011011001000111111) && ({row_reg, col_reg}<20'b00011011001001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00011011001001100110) && ({row_reg, col_reg}<20'b00011011001001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00011011001001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00011011001001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00011011001001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00011011001001101011) && ({row_reg, col_reg}<20'b00011011010100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00011011010100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00011011010100011111) && ({row_reg, col_reg}<20'b00011011010101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00011011010101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00011011010101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00011011010101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00011011010101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00011011010101010000) && ({row_reg, col_reg}<20'b00011011011000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00011011011000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00011011011000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00011011011000111000) && ({row_reg, col_reg}<20'b00011011011000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00011011011000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00011011011000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00011011011000111100) && ({row_reg, col_reg}<20'b00011011011000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00011011011000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00011011011000111111) && ({row_reg, col_reg}<20'b00011011011001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00011011011001100110) && ({row_reg, col_reg}<20'b00011011011001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00011011011001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00011011011001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00011011011001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00011011011001101011) && ({row_reg, col_reg}<20'b00011011100100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00011011100100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00011011100100011111) && ({row_reg, col_reg}<20'b00011011100101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00011011100101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00011011100101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00011011100101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00011011100101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00011011100101010000) && ({row_reg, col_reg}<20'b00011011101000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00011011101000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00011011101000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00011011101000111000) && ({row_reg, col_reg}<20'b00011011101000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00011011101000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00011011101000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00011011101000111100) && ({row_reg, col_reg}<20'b00011011101000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00011011101000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00011011101000111111) && ({row_reg, col_reg}<20'b00011011101001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00011011101001100110) && ({row_reg, col_reg}<20'b00011011101001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00011011101001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00011011101001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00011011101001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00011011101001101011) && ({row_reg, col_reg}<20'b00011011110100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00011011110100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00011011110100011111) && ({row_reg, col_reg}<20'b00011011110101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00011011110101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00011011110101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00011011110101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00011011110101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00011011110101010000) && ({row_reg, col_reg}<20'b00011011111000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00011011111000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00011011111000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00011011111000111000) && ({row_reg, col_reg}<20'b00011011111000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00011011111000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00011011111000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00011011111000111100) && ({row_reg, col_reg}<20'b00011011111000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00011011111000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00011011111000111111) && ({row_reg, col_reg}<20'b00011011111001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00011011111001100110) && ({row_reg, col_reg}<20'b00011011111001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00011011111001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00011011111001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00011011111001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00011011111001101011) && ({row_reg, col_reg}<20'b00011100000100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00011100000100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00011100000100011111) && ({row_reg, col_reg}<20'b00011100000101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00011100000101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00011100000101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00011100000101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00011100000101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00011100000101010000) && ({row_reg, col_reg}<20'b00011100001000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00011100001000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00011100001000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00011100001000111000) && ({row_reg, col_reg}<20'b00011100001000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00011100001000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00011100001000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00011100001000111100) && ({row_reg, col_reg}<20'b00011100001000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00011100001000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00011100001000111111) && ({row_reg, col_reg}<20'b00011100001001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00011100001001100110) && ({row_reg, col_reg}<20'b00011100001001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00011100001001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00011100001001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00011100001001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00011100001001101011) && ({row_reg, col_reg}<20'b00011100010100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00011100010100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00011100010100011111) && ({row_reg, col_reg}<20'b00011100010101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00011100010101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00011100010101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00011100010101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00011100010101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00011100010101010000) && ({row_reg, col_reg}<20'b00011100011000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00011100011000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00011100011000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00011100011000111000) && ({row_reg, col_reg}<20'b00011100011000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00011100011000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00011100011000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00011100011000111100) && ({row_reg, col_reg}<20'b00011100011000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00011100011000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00011100011000111111) && ({row_reg, col_reg}<20'b00011100011001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00011100011001100110) && ({row_reg, col_reg}<20'b00011100011001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00011100011001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00011100011001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00011100011001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00011100011001101011) && ({row_reg, col_reg}<20'b00011100100100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00011100100100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00011100100100011111) && ({row_reg, col_reg}<20'b00011100100101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00011100100101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00011100100101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00011100100101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00011100100101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00011100100101010000) && ({row_reg, col_reg}<20'b00011100101000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00011100101000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00011100101000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00011100101000111000) && ({row_reg, col_reg}<20'b00011100101000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00011100101000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00011100101000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00011100101000111100) && ({row_reg, col_reg}<20'b00011100101000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00011100101000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00011100101000111111) && ({row_reg, col_reg}<20'b00011100101001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00011100101001100110) && ({row_reg, col_reg}<20'b00011100101001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00011100101001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00011100101001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00011100101001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00011100101001101011) && ({row_reg, col_reg}<20'b00011100110100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00011100110100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00011100110100011111) && ({row_reg, col_reg}<20'b00011100110101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00011100110101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00011100110101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00011100110101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00011100110101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00011100110101010000) && ({row_reg, col_reg}<20'b00011100111000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00011100111000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00011100111000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00011100111000111000) && ({row_reg, col_reg}<20'b00011100111000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00011100111000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00011100111000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00011100111000111100) && ({row_reg, col_reg}<20'b00011100111000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00011100111000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00011100111000111111) && ({row_reg, col_reg}<20'b00011100111001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00011100111001100110) && ({row_reg, col_reg}<20'b00011100111001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00011100111001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00011100111001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00011100111001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00011100111001101011) && ({row_reg, col_reg}<20'b00011101000100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00011101000100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00011101000100011111) && ({row_reg, col_reg}<20'b00011101000101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00011101000101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00011101000101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00011101000101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00011101000101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00011101000101010000) && ({row_reg, col_reg}<20'b00011101001000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00011101001000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00011101001000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00011101001000111000) && ({row_reg, col_reg}<20'b00011101001000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00011101001000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00011101001000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00011101001000111100) && ({row_reg, col_reg}<20'b00011101001000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00011101001000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00011101001000111111) && ({row_reg, col_reg}<20'b00011101001001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00011101001001100110) && ({row_reg, col_reg}<20'b00011101001001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00011101001001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00011101001001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00011101001001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00011101001001101011) && ({row_reg, col_reg}<20'b00011101010100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00011101010100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00011101010100011111) && ({row_reg, col_reg}<20'b00011101010101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00011101010101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00011101010101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00011101010101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00011101010101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00011101010101010000) && ({row_reg, col_reg}<20'b00011101011000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00011101011000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00011101011000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00011101011000111000) && ({row_reg, col_reg}<20'b00011101011000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00011101011000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00011101011000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00011101011000111100) && ({row_reg, col_reg}<20'b00011101011000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00011101011000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00011101011000111111) && ({row_reg, col_reg}<20'b00011101011001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00011101011001100110) && ({row_reg, col_reg}<20'b00011101011001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00011101011001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00011101011001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00011101011001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00011101011001101011) && ({row_reg, col_reg}<20'b00011101100100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00011101100100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00011101100100011111) && ({row_reg, col_reg}<20'b00011101100101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00011101100101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00011101100101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00011101100101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00011101100101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00011101100101010000) && ({row_reg, col_reg}<20'b00011101101000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00011101101000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00011101101000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00011101101000111000) && ({row_reg, col_reg}<20'b00011101101000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00011101101000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00011101101000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00011101101000111100) && ({row_reg, col_reg}<20'b00011101101000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00011101101000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00011101101000111111) && ({row_reg, col_reg}<20'b00011101101001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00011101101001100110) && ({row_reg, col_reg}<20'b00011101101001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00011101101001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00011101101001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00011101101001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00011101101001101011) && ({row_reg, col_reg}<20'b00011101110100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00011101110100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00011101110100011111) && ({row_reg, col_reg}<20'b00011101110101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00011101110101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00011101110101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00011101110101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00011101110101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00011101110101010000) && ({row_reg, col_reg}<20'b00011101111000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00011101111000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00011101111000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00011101111000111000) && ({row_reg, col_reg}<20'b00011101111000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00011101111000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00011101111000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00011101111000111100) && ({row_reg, col_reg}<20'b00011101111000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00011101111000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00011101111000111111) && ({row_reg, col_reg}<20'b00011101111001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00011101111001100110) && ({row_reg, col_reg}<20'b00011101111001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00011101111001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00011101111001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00011101111001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00011101111001101011) && ({row_reg, col_reg}<20'b00011110000100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00011110000100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00011110000100011111) && ({row_reg, col_reg}<20'b00011110000101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00011110000101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00011110000101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00011110000101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00011110000101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00011110000101010000) && ({row_reg, col_reg}<20'b00011110001000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00011110001000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00011110001000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00011110001000111000) && ({row_reg, col_reg}<20'b00011110001000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00011110001000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00011110001000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00011110001000111100) && ({row_reg, col_reg}<20'b00011110001000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00011110001000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00011110001000111111) && ({row_reg, col_reg}<20'b00011110001001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00011110001001100110) && ({row_reg, col_reg}<20'b00011110001001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00011110001001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00011110001001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00011110001001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00011110001001101011) && ({row_reg, col_reg}<20'b00011110010100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00011110010100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00011110010100011111) && ({row_reg, col_reg}<20'b00011110010101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00011110010101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00011110010101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00011110010101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00011110010101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00011110010101010000) && ({row_reg, col_reg}<20'b00011110011000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00011110011000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00011110011000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00011110011000111000) && ({row_reg, col_reg}<20'b00011110011000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00011110011000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00011110011000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00011110011000111100) && ({row_reg, col_reg}<20'b00011110011000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00011110011000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00011110011000111111) && ({row_reg, col_reg}<20'b00011110011001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00011110011001100110) && ({row_reg, col_reg}<20'b00011110011001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00011110011001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00011110011001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00011110011001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00011110011001101011) && ({row_reg, col_reg}<20'b00011110100100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00011110100100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00011110100100011111) && ({row_reg, col_reg}<20'b00011110100101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00011110100101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00011110100101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00011110100101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00011110100101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00011110100101010000) && ({row_reg, col_reg}<20'b00011110101000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00011110101000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00011110101000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00011110101000111000) && ({row_reg, col_reg}<20'b00011110101000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00011110101000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00011110101000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00011110101000111100) && ({row_reg, col_reg}<20'b00011110101000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00011110101000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00011110101000111111) && ({row_reg, col_reg}<20'b00011110101001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00011110101001100110) && ({row_reg, col_reg}<20'b00011110101001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00011110101001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00011110101001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00011110101001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00011110101001101011) && ({row_reg, col_reg}<20'b00011110110100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00011110110100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00011110110100011111) && ({row_reg, col_reg}<20'b00011110110101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00011110110101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00011110110101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00011110110101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00011110110101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00011110110101010000) && ({row_reg, col_reg}<20'b00011110111000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00011110111000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00011110111000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00011110111000111000) && ({row_reg, col_reg}<20'b00011110111000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00011110111000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00011110111000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00011110111000111100) && ({row_reg, col_reg}<20'b00011110111000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00011110111000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00011110111000111111) && ({row_reg, col_reg}<20'b00011110111001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00011110111001100110) && ({row_reg, col_reg}<20'b00011110111001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00011110111001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00011110111001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00011110111001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00011110111001101011) && ({row_reg, col_reg}<20'b00011111000100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00011111000100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00011111000100011111) && ({row_reg, col_reg}<20'b00011111000101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00011111000101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00011111000101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00011111000101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00011111000101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00011111000101010000) && ({row_reg, col_reg}<20'b00011111001000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00011111001000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00011111001000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00011111001000111000) && ({row_reg, col_reg}<20'b00011111001000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00011111001000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00011111001000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00011111001000111100) && ({row_reg, col_reg}<20'b00011111001000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00011111001000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00011111001000111111) && ({row_reg, col_reg}<20'b00011111001001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00011111001001100110) && ({row_reg, col_reg}<20'b00011111001001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00011111001001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00011111001001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00011111001001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00011111001001101011) && ({row_reg, col_reg}<20'b00011111010100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00011111010100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00011111010100011111) && ({row_reg, col_reg}<20'b00011111010101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00011111010101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00011111010101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00011111010101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00011111010101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00011111010101010000) && ({row_reg, col_reg}<20'b00011111011000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00011111011000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00011111011000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00011111011000111000) && ({row_reg, col_reg}<20'b00011111011000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00011111011000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00011111011000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00011111011000111100) && ({row_reg, col_reg}<20'b00011111011000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00011111011000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00011111011000111111) && ({row_reg, col_reg}<20'b00011111011001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00011111011001100110) && ({row_reg, col_reg}<20'b00011111011001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00011111011001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00011111011001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00011111011001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00011111011001101011) && ({row_reg, col_reg}<20'b00011111100100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00011111100100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00011111100100011111) && ({row_reg, col_reg}<20'b00011111100101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00011111100101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00011111100101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00011111100101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00011111100101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00011111100101010000) && ({row_reg, col_reg}<20'b00011111101000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00011111101000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00011111101000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00011111101000111000) && ({row_reg, col_reg}<20'b00011111101000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00011111101000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00011111101000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00011111101000111100) && ({row_reg, col_reg}<20'b00011111101000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00011111101000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00011111101000111111) && ({row_reg, col_reg}<20'b00011111101001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00011111101001100110) && ({row_reg, col_reg}<20'b00011111101001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00011111101001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00011111101001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00011111101001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00011111101001101011) && ({row_reg, col_reg}<20'b00011111110100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00011111110100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00011111110100011111) && ({row_reg, col_reg}<20'b00011111110101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00011111110101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00011111110101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00011111110101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00011111110101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00011111110101010000) && ({row_reg, col_reg}<20'b00011111111000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00011111111000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00011111111000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00011111111000111000) && ({row_reg, col_reg}<20'b00011111111000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00011111111000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00011111111000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00011111111000111100) && ({row_reg, col_reg}<20'b00011111111000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00011111111000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00011111111000111111) && ({row_reg, col_reg}<20'b00011111111001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00011111111001100110) && ({row_reg, col_reg}<20'b00011111111001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00011111111001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00011111111001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00011111111001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00011111111001101011) && ({row_reg, col_reg}<20'b00100000000100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00100000000100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00100000000100011111) && ({row_reg, col_reg}<20'b00100000000101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00100000000101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00100000000101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00100000000101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00100000000101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00100000000101010000) && ({row_reg, col_reg}<20'b00100000001000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00100000001000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00100000001000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00100000001000111000) && ({row_reg, col_reg}<20'b00100000001000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00100000001000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00100000001000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00100000001000111100) && ({row_reg, col_reg}<20'b00100000001000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00100000001000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00100000001000111111) && ({row_reg, col_reg}<20'b00100000001001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00100000001001100110) && ({row_reg, col_reg}<20'b00100000001001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00100000001001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00100000001001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00100000001001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00100000001001101011) && ({row_reg, col_reg}<20'b00100000010100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00100000010100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00100000010100011111) && ({row_reg, col_reg}<20'b00100000010101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00100000010101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00100000010101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00100000010101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00100000010101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00100000010101010000) && ({row_reg, col_reg}<20'b00100000011000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00100000011000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00100000011000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00100000011000111000) && ({row_reg, col_reg}<20'b00100000011000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00100000011000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00100000011000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00100000011000111100) && ({row_reg, col_reg}<20'b00100000011000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00100000011000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00100000011000111111) && ({row_reg, col_reg}<20'b00100000011001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00100000011001100110) && ({row_reg, col_reg}<20'b00100000011001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00100000011001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00100000011001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00100000011001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00100000011001101011) && ({row_reg, col_reg}<20'b00100000100100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00100000100100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00100000100100011111) && ({row_reg, col_reg}<20'b00100000100101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00100000100101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00100000100101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00100000100101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00100000100101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00100000100101010000) && ({row_reg, col_reg}<20'b00100000101000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00100000101000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00100000101000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00100000101000111000) && ({row_reg, col_reg}<20'b00100000101000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00100000101000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00100000101000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00100000101000111100) && ({row_reg, col_reg}<20'b00100000101000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00100000101000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00100000101000111111) && ({row_reg, col_reg}<20'b00100000101001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00100000101001100110) && ({row_reg, col_reg}<20'b00100000101001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00100000101001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00100000101001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00100000101001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00100000101001101011) && ({row_reg, col_reg}<20'b00100000110100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00100000110100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00100000110100011111) && ({row_reg, col_reg}<20'b00100000110101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00100000110101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00100000110101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00100000110101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00100000110101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00100000110101010000) && ({row_reg, col_reg}<20'b00100000111000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00100000111000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00100000111000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00100000111000111000) && ({row_reg, col_reg}<20'b00100000111000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00100000111000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00100000111000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00100000111000111100) && ({row_reg, col_reg}<20'b00100000111000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00100000111000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00100000111000111111) && ({row_reg, col_reg}<20'b00100000111001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00100000111001100110) && ({row_reg, col_reg}<20'b00100000111001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00100000111001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00100000111001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00100000111001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00100000111001101011) && ({row_reg, col_reg}<20'b00100001000100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00100001000100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00100001000100011111) && ({row_reg, col_reg}<20'b00100001000101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00100001000101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00100001000101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00100001000101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00100001000101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00100001000101010000) && ({row_reg, col_reg}<20'b00100001001000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00100001001000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00100001001000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00100001001000111000) && ({row_reg, col_reg}<20'b00100001001000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00100001001000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00100001001000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00100001001000111100) && ({row_reg, col_reg}<20'b00100001001000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00100001001000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00100001001000111111) && ({row_reg, col_reg}<20'b00100001001001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00100001001001100110) && ({row_reg, col_reg}<20'b00100001001001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00100001001001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00100001001001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00100001001001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00100001001001101011) && ({row_reg, col_reg}<20'b00100001010100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00100001010100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00100001010100011111) && ({row_reg, col_reg}<20'b00100001010101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00100001010101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00100001010101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00100001010101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00100001010101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00100001010101010000) && ({row_reg, col_reg}<20'b00100001011000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00100001011000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00100001011000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00100001011000111000) && ({row_reg, col_reg}<20'b00100001011000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00100001011000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00100001011000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00100001011000111100) && ({row_reg, col_reg}<20'b00100001011000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00100001011000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00100001011000111111) && ({row_reg, col_reg}<20'b00100001011001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00100001011001100110) && ({row_reg, col_reg}<20'b00100001011001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00100001011001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00100001011001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00100001011001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00100001011001101011) && ({row_reg, col_reg}<20'b00100001100100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00100001100100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00100001100100011111) && ({row_reg, col_reg}<20'b00100001100101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00100001100101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00100001100101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00100001100101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00100001100101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00100001100101010000) && ({row_reg, col_reg}<20'b00100001101000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00100001101000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00100001101000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00100001101000111000) && ({row_reg, col_reg}<20'b00100001101000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00100001101000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00100001101000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00100001101000111100) && ({row_reg, col_reg}<20'b00100001101000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00100001101000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00100001101000111111) && ({row_reg, col_reg}<20'b00100001101001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00100001101001100110) && ({row_reg, col_reg}<20'b00100001101001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00100001101001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00100001101001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00100001101001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00100001101001101011) && ({row_reg, col_reg}<20'b00100001110100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00100001110100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00100001110100011111) && ({row_reg, col_reg}<20'b00100001110101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00100001110101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00100001110101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00100001110101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00100001110101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00100001110101010000) && ({row_reg, col_reg}<20'b00100001111000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00100001111000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00100001111000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00100001111000111000) && ({row_reg, col_reg}<20'b00100001111000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00100001111000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00100001111000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00100001111000111100) && ({row_reg, col_reg}<20'b00100001111000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00100001111000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00100001111000111111) && ({row_reg, col_reg}<20'b00100001111001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00100001111001100110) && ({row_reg, col_reg}<20'b00100001111001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00100001111001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00100001111001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00100001111001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00100001111001101011) && ({row_reg, col_reg}<20'b00100010000100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00100010000100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00100010000100011111) && ({row_reg, col_reg}<20'b00100010000101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00100010000101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00100010000101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00100010000101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00100010000101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00100010000101010000) && ({row_reg, col_reg}<20'b00100010001000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00100010001000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00100010001000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00100010001000111000) && ({row_reg, col_reg}<20'b00100010001000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00100010001000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00100010001000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00100010001000111100) && ({row_reg, col_reg}<20'b00100010001000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00100010001000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00100010001000111111) && ({row_reg, col_reg}<20'b00100010001001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00100010001001100110) && ({row_reg, col_reg}<20'b00100010001001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00100010001001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00100010001001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00100010001001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00100010001001101011) && ({row_reg, col_reg}<20'b00100010010100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00100010010100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00100010010100011111) && ({row_reg, col_reg}<20'b00100010010101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00100010010101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00100010010101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00100010010101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00100010010101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00100010010101010000) && ({row_reg, col_reg}<20'b00100010011000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00100010011000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00100010011000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00100010011000111000) && ({row_reg, col_reg}<20'b00100010011000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00100010011000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00100010011000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00100010011000111100) && ({row_reg, col_reg}<20'b00100010011000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00100010011000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00100010011000111111) && ({row_reg, col_reg}<20'b00100010011001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00100010011001100110) && ({row_reg, col_reg}<20'b00100010011001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00100010011001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00100010011001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00100010011001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00100010011001101011) && ({row_reg, col_reg}<20'b00100010100100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00100010100100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00100010100100011111) && ({row_reg, col_reg}<20'b00100010100101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00100010100101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00100010100101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00100010100101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00100010100101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00100010100101010000) && ({row_reg, col_reg}<20'b00100010101000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00100010101000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00100010101000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00100010101000111000) && ({row_reg, col_reg}<20'b00100010101000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00100010101000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00100010101000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00100010101000111100) && ({row_reg, col_reg}<20'b00100010101000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00100010101000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00100010101000111111) && ({row_reg, col_reg}<20'b00100010101001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00100010101001100110) && ({row_reg, col_reg}<20'b00100010101001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00100010101001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00100010101001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00100010101001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00100010101001101011) && ({row_reg, col_reg}<20'b00100010110100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00100010110100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00100010110100011111) && ({row_reg, col_reg}<20'b00100010110101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00100010110101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00100010110101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00100010110101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00100010110101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00100010110101010000) && ({row_reg, col_reg}<20'b00100010111000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00100010111000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00100010111000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00100010111000111000) && ({row_reg, col_reg}<20'b00100010111000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00100010111000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00100010111000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00100010111000111100) && ({row_reg, col_reg}<20'b00100010111000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00100010111000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00100010111000111111) && ({row_reg, col_reg}<20'b00100010111001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00100010111001100110) && ({row_reg, col_reg}<20'b00100010111001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00100010111001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00100010111001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00100010111001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00100010111001101011) && ({row_reg, col_reg}<20'b00100011000100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00100011000100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00100011000100011111) && ({row_reg, col_reg}<20'b00100011000101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00100011000101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00100011000101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00100011000101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00100011000101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00100011000101010000) && ({row_reg, col_reg}<20'b00100011001000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00100011001000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00100011001000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00100011001000111000) && ({row_reg, col_reg}<20'b00100011001000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00100011001000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00100011001000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00100011001000111100) && ({row_reg, col_reg}<20'b00100011001000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00100011001000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00100011001000111111) && ({row_reg, col_reg}<20'b00100011001001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00100011001001100110) && ({row_reg, col_reg}<20'b00100011001001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00100011001001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00100011001001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00100011001001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00100011001001101011) && ({row_reg, col_reg}<20'b00100011010100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00100011010100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00100011010100011111) && ({row_reg, col_reg}<20'b00100011010101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00100011010101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00100011010101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00100011010101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00100011010101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00100011010101010000) && ({row_reg, col_reg}<20'b00100011011000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00100011011000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00100011011000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00100011011000111000) && ({row_reg, col_reg}<20'b00100011011000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00100011011000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00100011011000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00100011011000111100) && ({row_reg, col_reg}<20'b00100011011000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00100011011000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00100011011000111111) && ({row_reg, col_reg}<20'b00100011011001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00100011011001100110) && ({row_reg, col_reg}<20'b00100011011001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00100011011001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00100011011001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00100011011001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00100011011001101011) && ({row_reg, col_reg}<20'b00100011100100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00100011100100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00100011100100011111) && ({row_reg, col_reg}<20'b00100011100101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00100011100101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00100011100101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00100011100101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00100011100101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00100011100101010000) && ({row_reg, col_reg}<20'b00100011101000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00100011101000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00100011101000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00100011101000111000) && ({row_reg, col_reg}<20'b00100011101000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00100011101000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00100011101000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00100011101000111100) && ({row_reg, col_reg}<20'b00100011101000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00100011101000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00100011101000111111) && ({row_reg, col_reg}<20'b00100011101001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00100011101001100110) && ({row_reg, col_reg}<20'b00100011101001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00100011101001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00100011101001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00100011101001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00100011101001101011) && ({row_reg, col_reg}<20'b00100011110100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00100011110100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00100011110100011111) && ({row_reg, col_reg}<20'b00100011110101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00100011110101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00100011110101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00100011110101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00100011110101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00100011110101010000) && ({row_reg, col_reg}<20'b00100011111000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00100011111000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00100011111000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00100011111000111000) && ({row_reg, col_reg}<20'b00100011111000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00100011111000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00100011111000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00100011111000111100) && ({row_reg, col_reg}<20'b00100011111000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00100011111000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00100011111000111111) && ({row_reg, col_reg}<20'b00100011111001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00100011111001100110) && ({row_reg, col_reg}<20'b00100011111001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00100011111001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00100011111001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00100011111001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00100011111001101011) && ({row_reg, col_reg}<20'b00100100000100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00100100000100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00100100000100011111) && ({row_reg, col_reg}<20'b00100100000101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00100100000101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00100100000101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00100100000101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00100100000101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00100100000101010000) && ({row_reg, col_reg}<20'b00100100001000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00100100001000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00100100001000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00100100001000111000) && ({row_reg, col_reg}<20'b00100100001000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00100100001000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00100100001000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00100100001000111100) && ({row_reg, col_reg}<20'b00100100001000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00100100001000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00100100001000111111) && ({row_reg, col_reg}<20'b00100100001001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00100100001001100110) && ({row_reg, col_reg}<20'b00100100001001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00100100001001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00100100001001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00100100001001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00100100001001101011) && ({row_reg, col_reg}<20'b00100100010100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00100100010100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00100100010100011111) && ({row_reg, col_reg}<20'b00100100010101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00100100010101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00100100010101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00100100010101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00100100010101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00100100010101010000) && ({row_reg, col_reg}<20'b00100100011000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00100100011000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00100100011000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00100100011000111000) && ({row_reg, col_reg}<20'b00100100011000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00100100011000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00100100011000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00100100011000111100) && ({row_reg, col_reg}<20'b00100100011000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00100100011000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00100100011000111111) && ({row_reg, col_reg}<20'b00100100011001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00100100011001100110) && ({row_reg, col_reg}<20'b00100100011001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00100100011001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00100100011001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00100100011001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00100100011001101011) && ({row_reg, col_reg}<20'b00100100100100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00100100100100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00100100100100011111) && ({row_reg, col_reg}<20'b00100100100101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00100100100101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00100100100101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00100100100101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00100100100101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00100100100101010000) && ({row_reg, col_reg}<20'b00100100101000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00100100101000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00100100101000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00100100101000111000) && ({row_reg, col_reg}<20'b00100100101000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00100100101000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00100100101000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00100100101000111100) && ({row_reg, col_reg}<20'b00100100101000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00100100101000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00100100101000111111) && ({row_reg, col_reg}<20'b00100100101001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00100100101001100110) && ({row_reg, col_reg}<20'b00100100101001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00100100101001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00100100101001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00100100101001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00100100101001101011) && ({row_reg, col_reg}<20'b00100100110100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00100100110100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00100100110100011111) && ({row_reg, col_reg}<20'b00100100110101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00100100110101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00100100110101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00100100110101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00100100110101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00100100110101010000) && ({row_reg, col_reg}<20'b00100100111000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00100100111000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00100100111000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00100100111000111000) && ({row_reg, col_reg}<20'b00100100111000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00100100111000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00100100111000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00100100111000111100) && ({row_reg, col_reg}<20'b00100100111000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00100100111000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00100100111000111111) && ({row_reg, col_reg}<20'b00100100111001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00100100111001100110) && ({row_reg, col_reg}<20'b00100100111001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00100100111001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00100100111001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00100100111001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00100100111001101011) && ({row_reg, col_reg}<20'b00100101000100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00100101000100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00100101000100011111) && ({row_reg, col_reg}<20'b00100101000101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00100101000101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00100101000101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00100101000101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00100101000101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00100101000101010000) && ({row_reg, col_reg}<20'b00100101001000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00100101001000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00100101001000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00100101001000111000) && ({row_reg, col_reg}<20'b00100101001000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00100101001000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00100101001000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00100101001000111100) && ({row_reg, col_reg}<20'b00100101001000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00100101001000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00100101001000111111) && ({row_reg, col_reg}<20'b00100101001001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00100101001001100110) && ({row_reg, col_reg}<20'b00100101001001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00100101001001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00100101001001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00100101001001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00100101001001101011) && ({row_reg, col_reg}<20'b00100101010100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00100101010100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00100101010100011111) && ({row_reg, col_reg}<20'b00100101010101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00100101010101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00100101010101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00100101010101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00100101010101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00100101010101010000) && ({row_reg, col_reg}<20'b00100101011000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00100101011000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00100101011000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00100101011000111000) && ({row_reg, col_reg}<20'b00100101011000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00100101011000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00100101011000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00100101011000111100) && ({row_reg, col_reg}<20'b00100101011000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00100101011000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00100101011000111111) && ({row_reg, col_reg}<20'b00100101011001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00100101011001100110) && ({row_reg, col_reg}<20'b00100101011001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00100101011001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00100101011001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00100101011001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00100101011001101011) && ({row_reg, col_reg}<20'b00100101100100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00100101100100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00100101100100011111) && ({row_reg, col_reg}<20'b00100101100101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00100101100101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00100101100101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00100101100101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00100101100101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00100101100101010000) && ({row_reg, col_reg}<20'b00100101101000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00100101101000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00100101101000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00100101101000111000) && ({row_reg, col_reg}<20'b00100101101000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00100101101000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00100101101000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00100101101000111100) && ({row_reg, col_reg}<20'b00100101101000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00100101101000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00100101101000111111) && ({row_reg, col_reg}<20'b00100101101001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00100101101001100110) && ({row_reg, col_reg}<20'b00100101101001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00100101101001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00100101101001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00100101101001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00100101101001101011) && ({row_reg, col_reg}<20'b00100101110100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00100101110100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00100101110100011111) && ({row_reg, col_reg}<20'b00100101110101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00100101110101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00100101110101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00100101110101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00100101110101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00100101110101010000) && ({row_reg, col_reg}<20'b00100101111000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00100101111000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00100101111000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00100101111000111000) && ({row_reg, col_reg}<20'b00100101111000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00100101111000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00100101111000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00100101111000111100) && ({row_reg, col_reg}<20'b00100101111000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00100101111000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00100101111000111111) && ({row_reg, col_reg}<20'b00100101111001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00100101111001100110) && ({row_reg, col_reg}<20'b00100101111001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00100101111001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00100101111001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00100101111001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00100101111001101011) && ({row_reg, col_reg}<20'b00100110000100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00100110000100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00100110000100011111) && ({row_reg, col_reg}<20'b00100110000101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00100110000101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00100110000101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00100110000101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00100110000101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00100110000101010000) && ({row_reg, col_reg}<20'b00100110001000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00100110001000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00100110001000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00100110001000111000) && ({row_reg, col_reg}<20'b00100110001000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00100110001000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00100110001000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00100110001000111100) && ({row_reg, col_reg}<20'b00100110001000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00100110001000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00100110001000111111) && ({row_reg, col_reg}<20'b00100110001001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00100110001001100110) && ({row_reg, col_reg}<20'b00100110001001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00100110001001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00100110001001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00100110001001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00100110001001101011) && ({row_reg, col_reg}<20'b00100110010100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00100110010100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00100110010100011111) && ({row_reg, col_reg}<20'b00100110010101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00100110010101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00100110010101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00100110010101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00100110010101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00100110010101010000) && ({row_reg, col_reg}<20'b00100110011000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00100110011000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00100110011000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00100110011000111000) && ({row_reg, col_reg}<20'b00100110011000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00100110011000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00100110011000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00100110011000111100) && ({row_reg, col_reg}<20'b00100110011000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00100110011000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00100110011000111111) && ({row_reg, col_reg}<20'b00100110011001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00100110011001100110) && ({row_reg, col_reg}<20'b00100110011001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00100110011001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00100110011001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00100110011001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00100110011001101011) && ({row_reg, col_reg}<20'b00100110100100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00100110100100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00100110100100011111) && ({row_reg, col_reg}<20'b00100110100101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00100110100101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00100110100101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00100110100101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00100110100101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00100110100101010000) && ({row_reg, col_reg}<20'b00100110101000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00100110101000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00100110101000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00100110101000111000) && ({row_reg, col_reg}<20'b00100110101000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00100110101000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00100110101000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00100110101000111100) && ({row_reg, col_reg}<20'b00100110101000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00100110101000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00100110101000111111) && ({row_reg, col_reg}<20'b00100110101001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00100110101001100110) && ({row_reg, col_reg}<20'b00100110101001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00100110101001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00100110101001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00100110101001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00100110101001101011) && ({row_reg, col_reg}<20'b00100110110100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00100110110100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00100110110100011111) && ({row_reg, col_reg}<20'b00100110110101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00100110110101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00100110110101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00100110110101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00100110110101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00100110110101010000) && ({row_reg, col_reg}<20'b00100110111000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00100110111000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00100110111000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00100110111000111000) && ({row_reg, col_reg}<20'b00100110111000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00100110111000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00100110111000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00100110111000111100) && ({row_reg, col_reg}<20'b00100110111000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00100110111000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00100110111000111111) && ({row_reg, col_reg}<20'b00100110111001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00100110111001100110) && ({row_reg, col_reg}<20'b00100110111001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00100110111001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00100110111001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00100110111001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00100110111001101011) && ({row_reg, col_reg}<20'b00100111000100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00100111000100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00100111000100011111) && ({row_reg, col_reg}<20'b00100111000101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00100111000101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00100111000101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00100111000101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00100111000101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00100111000101010000) && ({row_reg, col_reg}<20'b00100111001000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00100111001000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00100111001000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00100111001000111000) && ({row_reg, col_reg}<20'b00100111001000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00100111001000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00100111001000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00100111001000111100) && ({row_reg, col_reg}<20'b00100111001000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00100111001000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00100111001000111111) && ({row_reg, col_reg}<20'b00100111001001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00100111001001100110) && ({row_reg, col_reg}<20'b00100111001001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00100111001001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00100111001001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00100111001001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00100111001001101011) && ({row_reg, col_reg}<20'b00100111010100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00100111010100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00100111010100011111) && ({row_reg, col_reg}<20'b00100111010101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00100111010101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00100111010101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00100111010101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00100111010101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00100111010101010000) && ({row_reg, col_reg}<20'b00100111011000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00100111011000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00100111011000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00100111011000111000) && ({row_reg, col_reg}<20'b00100111011000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00100111011000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00100111011000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00100111011000111100) && ({row_reg, col_reg}<20'b00100111011000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00100111011000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00100111011000111111) && ({row_reg, col_reg}<20'b00100111011001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00100111011001100110) && ({row_reg, col_reg}<20'b00100111011001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00100111011001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00100111011001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00100111011001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00100111011001101011) && ({row_reg, col_reg}<20'b00100111100100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00100111100100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00100111100100011111) && ({row_reg, col_reg}<20'b00100111100101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00100111100101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00100111100101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00100111100101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00100111100101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00100111100101010000) && ({row_reg, col_reg}<20'b00100111101000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00100111101000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00100111101000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00100111101000111000) && ({row_reg, col_reg}<20'b00100111101000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00100111101000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00100111101000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00100111101000111100) && ({row_reg, col_reg}<20'b00100111101000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00100111101000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00100111101000111111) && ({row_reg, col_reg}<20'b00100111101001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00100111101001100110) && ({row_reg, col_reg}<20'b00100111101001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00100111101001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00100111101001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00100111101001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00100111101001101011) && ({row_reg, col_reg}<20'b00100111110100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00100111110100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00100111110100011111) && ({row_reg, col_reg}<20'b00100111110101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00100111110101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00100111110101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00100111110101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00100111110101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00100111110101010000) && ({row_reg, col_reg}<20'b00100111111000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00100111111000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00100111111000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00100111111000111000) && ({row_reg, col_reg}<20'b00100111111000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00100111111000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00100111111000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00100111111000111100) && ({row_reg, col_reg}<20'b00100111111000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00100111111000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00100111111000111111) && ({row_reg, col_reg}<20'b00100111111001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00100111111001100110) && ({row_reg, col_reg}<20'b00100111111001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00100111111001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00100111111001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00100111111001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00100111111001101011) && ({row_reg, col_reg}<20'b00101000000100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00101000000100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00101000000100011111) && ({row_reg, col_reg}<20'b00101000000101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00101000000101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00101000000101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00101000000101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00101000000101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00101000000101010000) && ({row_reg, col_reg}<20'b00101000001000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00101000001000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00101000001000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00101000001000111000) && ({row_reg, col_reg}<20'b00101000001000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00101000001000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00101000001000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00101000001000111100) && ({row_reg, col_reg}<20'b00101000001000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00101000001000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00101000001000111111) && ({row_reg, col_reg}<20'b00101000001001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00101000001001100110) && ({row_reg, col_reg}<20'b00101000001001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00101000001001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00101000001001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00101000001001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00101000001001101011) && ({row_reg, col_reg}<20'b00101000010100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00101000010100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00101000010100011111) && ({row_reg, col_reg}<20'b00101000010101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00101000010101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00101000010101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00101000010101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00101000010101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00101000010101010000) && ({row_reg, col_reg}<20'b00101000011000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00101000011000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00101000011000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00101000011000111000) && ({row_reg, col_reg}<20'b00101000011000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00101000011000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00101000011000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00101000011000111100) && ({row_reg, col_reg}<20'b00101000011000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00101000011000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00101000011000111111) && ({row_reg, col_reg}<20'b00101000011001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00101000011001100110) && ({row_reg, col_reg}<20'b00101000011001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00101000011001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00101000011001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00101000011001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00101000011001101011) && ({row_reg, col_reg}<20'b00101000100100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00101000100100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00101000100100011111) && ({row_reg, col_reg}<20'b00101000100101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00101000100101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00101000100101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00101000100101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00101000100101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00101000100101010000) && ({row_reg, col_reg}<20'b00101000101000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00101000101000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00101000101000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00101000101000111000) && ({row_reg, col_reg}<20'b00101000101000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00101000101000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00101000101000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00101000101000111100) && ({row_reg, col_reg}<20'b00101000101000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00101000101000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00101000101000111111) && ({row_reg, col_reg}<20'b00101000101001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00101000101001100110) && ({row_reg, col_reg}<20'b00101000101001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00101000101001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00101000101001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00101000101001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00101000101001101011) && ({row_reg, col_reg}<20'b00101000110100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00101000110100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00101000110100011111) && ({row_reg, col_reg}<20'b00101000110101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00101000110101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00101000110101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00101000110101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00101000110101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00101000110101010000) && ({row_reg, col_reg}<20'b00101000111000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00101000111000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00101000111000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00101000111000111000) && ({row_reg, col_reg}<20'b00101000111000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00101000111000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00101000111000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00101000111000111100) && ({row_reg, col_reg}<20'b00101000111000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00101000111000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00101000111000111111) && ({row_reg, col_reg}<20'b00101000111001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00101000111001100110) && ({row_reg, col_reg}<20'b00101000111001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00101000111001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00101000111001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00101000111001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00101000111001101011) && ({row_reg, col_reg}<20'b00101001000100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00101001000100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00101001000100011111) && ({row_reg, col_reg}<20'b00101001000101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00101001000101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00101001000101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00101001000101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00101001000101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00101001000101010000) && ({row_reg, col_reg}<20'b00101001001000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00101001001000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00101001001000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00101001001000111000) && ({row_reg, col_reg}<20'b00101001001000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00101001001000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00101001001000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00101001001000111100) && ({row_reg, col_reg}<20'b00101001001000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00101001001000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00101001001000111111) && ({row_reg, col_reg}<20'b00101001001001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00101001001001100110) && ({row_reg, col_reg}<20'b00101001001001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00101001001001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00101001001001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00101001001001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00101001001001101011) && ({row_reg, col_reg}<20'b00101001010100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00101001010100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00101001010100011111) && ({row_reg, col_reg}<20'b00101001010101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00101001010101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00101001010101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00101001010101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00101001010101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00101001010101010000) && ({row_reg, col_reg}<20'b00101001011000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00101001011000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00101001011000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00101001011000111000) && ({row_reg, col_reg}<20'b00101001011000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00101001011000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00101001011000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00101001011000111100) && ({row_reg, col_reg}<20'b00101001011000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00101001011000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00101001011000111111) && ({row_reg, col_reg}<20'b00101001011001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00101001011001100110) && ({row_reg, col_reg}<20'b00101001011001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00101001011001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00101001011001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00101001011001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00101001011001101011) && ({row_reg, col_reg}<20'b00101001100100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00101001100100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00101001100100011111) && ({row_reg, col_reg}<20'b00101001100101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00101001100101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00101001100101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00101001100101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00101001100101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00101001100101010000) && ({row_reg, col_reg}<20'b00101001101000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00101001101000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00101001101000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00101001101000111000) && ({row_reg, col_reg}<20'b00101001101000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00101001101000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00101001101000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00101001101000111100) && ({row_reg, col_reg}<20'b00101001101000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00101001101000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00101001101000111111) && ({row_reg, col_reg}<20'b00101001101001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00101001101001100110) && ({row_reg, col_reg}<20'b00101001101001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00101001101001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00101001101001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00101001101001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00101001101001101011) && ({row_reg, col_reg}<20'b00101001110100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00101001110100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00101001110100011111) && ({row_reg, col_reg}<20'b00101001110101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00101001110101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00101001110101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00101001110101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00101001110101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00101001110101010000) && ({row_reg, col_reg}<20'b00101001111000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00101001111000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00101001111000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00101001111000111000) && ({row_reg, col_reg}<20'b00101001111000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00101001111000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00101001111000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00101001111000111100) && ({row_reg, col_reg}<20'b00101001111000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00101001111000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00101001111000111111) && ({row_reg, col_reg}<20'b00101001111001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00101001111001100110) && ({row_reg, col_reg}<20'b00101001111001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00101001111001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00101001111001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00101001111001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00101001111001101011) && ({row_reg, col_reg}<20'b00101010000100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00101010000100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00101010000100011111) && ({row_reg, col_reg}<20'b00101010000101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00101010000101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00101010000101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00101010000101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00101010000101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00101010000101010000) && ({row_reg, col_reg}<20'b00101010001000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00101010001000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00101010001000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00101010001000111000) && ({row_reg, col_reg}<20'b00101010001000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00101010001000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00101010001000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00101010001000111100) && ({row_reg, col_reg}<20'b00101010001000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00101010001000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00101010001000111111) && ({row_reg, col_reg}<20'b00101010001001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00101010001001100110) && ({row_reg, col_reg}<20'b00101010001001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00101010001001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00101010001001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00101010001001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00101010001001101011) && ({row_reg, col_reg}<20'b00101010010100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00101010010100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00101010010100011111) && ({row_reg, col_reg}<20'b00101010010101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00101010010101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00101010010101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00101010010101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00101010010101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00101010010101010000) && ({row_reg, col_reg}<20'b00101010011000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00101010011000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00101010011000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00101010011000111000) && ({row_reg, col_reg}<20'b00101010011000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00101010011000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00101010011000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00101010011000111100) && ({row_reg, col_reg}<20'b00101010011000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00101010011000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00101010011000111111) && ({row_reg, col_reg}<20'b00101010011001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00101010011001100110) && ({row_reg, col_reg}<20'b00101010011001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00101010011001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00101010011001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00101010011001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00101010011001101011) && ({row_reg, col_reg}<20'b00101010100100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00101010100100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00101010100100011111) && ({row_reg, col_reg}<20'b00101010100101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00101010100101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00101010100101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00101010100101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00101010100101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00101010100101010000) && ({row_reg, col_reg}<20'b00101010101000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00101010101000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00101010101000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00101010101000111000) && ({row_reg, col_reg}<20'b00101010101000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00101010101000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00101010101000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00101010101000111100) && ({row_reg, col_reg}<20'b00101010101000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00101010101000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00101010101000111111) && ({row_reg, col_reg}<20'b00101010101001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00101010101001100110) && ({row_reg, col_reg}<20'b00101010101001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00101010101001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00101010101001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00101010101001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00101010101001101011) && ({row_reg, col_reg}<20'b00101010110100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00101010110100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00101010110100011111) && ({row_reg, col_reg}<20'b00101010110101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00101010110101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00101010110101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00101010110101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00101010110101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00101010110101010000) && ({row_reg, col_reg}<20'b00101010111000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00101010111000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00101010111000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00101010111000111000) && ({row_reg, col_reg}<20'b00101010111000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00101010111000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00101010111000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00101010111000111100) && ({row_reg, col_reg}<20'b00101010111000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00101010111000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00101010111000111111) && ({row_reg, col_reg}<20'b00101010111001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00101010111001100110) && ({row_reg, col_reg}<20'b00101010111001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00101010111001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00101010111001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00101010111001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00101010111001101011) && ({row_reg, col_reg}<20'b00101011000100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00101011000100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00101011000100011111) && ({row_reg, col_reg}<20'b00101011000101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00101011000101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00101011000101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00101011000101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00101011000101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00101011000101010000) && ({row_reg, col_reg}<20'b00101011001000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00101011001000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00101011001000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00101011001000111000) && ({row_reg, col_reg}<20'b00101011001000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00101011001000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00101011001000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00101011001000111100) && ({row_reg, col_reg}<20'b00101011001000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00101011001000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00101011001000111111) && ({row_reg, col_reg}<20'b00101011001001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00101011001001100110) && ({row_reg, col_reg}<20'b00101011001001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00101011001001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00101011001001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00101011001001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00101011001001101011) && ({row_reg, col_reg}<20'b00101011010100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00101011010100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00101011010100011111) && ({row_reg, col_reg}<20'b00101011010101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00101011010101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00101011010101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00101011010101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00101011010101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00101011010101010000) && ({row_reg, col_reg}<20'b00101011011000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00101011011000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00101011011000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00101011011000111000) && ({row_reg, col_reg}<20'b00101011011000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00101011011000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00101011011000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00101011011000111100) && ({row_reg, col_reg}<20'b00101011011000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00101011011000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00101011011000111111) && ({row_reg, col_reg}<20'b00101011011001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00101011011001100110) && ({row_reg, col_reg}<20'b00101011011001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00101011011001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00101011011001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00101011011001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00101011011001101011) && ({row_reg, col_reg}<20'b00101011100100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00101011100100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00101011100100011111) && ({row_reg, col_reg}<20'b00101011100101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00101011100101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00101011100101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00101011100101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00101011100101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00101011100101010000) && ({row_reg, col_reg}<20'b00101011101000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00101011101000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00101011101000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00101011101000111000) && ({row_reg, col_reg}<20'b00101011101000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00101011101000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00101011101000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00101011101000111100) && ({row_reg, col_reg}<20'b00101011101000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00101011101000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00101011101000111111) && ({row_reg, col_reg}<20'b00101011101001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00101011101001100110) && ({row_reg, col_reg}<20'b00101011101001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00101011101001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00101011101001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00101011101001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00101011101001101011) && ({row_reg, col_reg}<20'b00101011110100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00101011110100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00101011110100011111) && ({row_reg, col_reg}<20'b00101011110101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00101011110101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00101011110101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00101011110101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00101011110101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00101011110101010000) && ({row_reg, col_reg}<20'b00101011111000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00101011111000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00101011111000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00101011111000111000) && ({row_reg, col_reg}<20'b00101011111000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00101011111000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00101011111000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00101011111000111100) && ({row_reg, col_reg}<20'b00101011111000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00101011111000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00101011111000111111) && ({row_reg, col_reg}<20'b00101011111001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00101011111001100110) && ({row_reg, col_reg}<20'b00101011111001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00101011111001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00101011111001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00101011111001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00101011111001101011) && ({row_reg, col_reg}<20'b00101100000100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00101100000100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00101100000100011111) && ({row_reg, col_reg}<20'b00101100000101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00101100000101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00101100000101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00101100000101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00101100000101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00101100000101010000) && ({row_reg, col_reg}<20'b00101100001000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00101100001000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00101100001000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00101100001000111000) && ({row_reg, col_reg}<20'b00101100001000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00101100001000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00101100001000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00101100001000111100) && ({row_reg, col_reg}<20'b00101100001000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00101100001000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00101100001000111111) && ({row_reg, col_reg}<20'b00101100001001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00101100001001100110) && ({row_reg, col_reg}<20'b00101100001001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00101100001001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00101100001001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00101100001001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00101100001001101011) && ({row_reg, col_reg}<20'b00101100010100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00101100010100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00101100010100011111) && ({row_reg, col_reg}<20'b00101100010101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00101100010101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00101100010101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00101100010101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00101100010101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00101100010101010000) && ({row_reg, col_reg}<20'b00101100011000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00101100011000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00101100011000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00101100011000111000) && ({row_reg, col_reg}<20'b00101100011000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00101100011000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00101100011000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00101100011000111100) && ({row_reg, col_reg}<20'b00101100011000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00101100011000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00101100011000111111) && ({row_reg, col_reg}<20'b00101100011001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00101100011001100110) && ({row_reg, col_reg}<20'b00101100011001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00101100011001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00101100011001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00101100011001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00101100011001101011) && ({row_reg, col_reg}<20'b00101100100100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00101100100100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00101100100100011111) && ({row_reg, col_reg}<20'b00101100100101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00101100100101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00101100100101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00101100100101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00101100100101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00101100100101010000) && ({row_reg, col_reg}<20'b00101100101000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00101100101000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00101100101000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00101100101000111000) && ({row_reg, col_reg}<20'b00101100101000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00101100101000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00101100101000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00101100101000111100) && ({row_reg, col_reg}<20'b00101100101000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00101100101000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00101100101000111111) && ({row_reg, col_reg}<20'b00101100101001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00101100101001100110) && ({row_reg, col_reg}<20'b00101100101001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00101100101001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00101100101001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00101100101001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00101100101001101011) && ({row_reg, col_reg}<20'b00101100110100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00101100110100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00101100110100011111) && ({row_reg, col_reg}<20'b00101100110101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00101100110101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00101100110101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00101100110101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00101100110101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00101100110101010000) && ({row_reg, col_reg}<20'b00101100111000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00101100111000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00101100111000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00101100111000111000) && ({row_reg, col_reg}<20'b00101100111000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00101100111000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00101100111000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00101100111000111100) && ({row_reg, col_reg}<20'b00101100111000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00101100111000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00101100111000111111) && ({row_reg, col_reg}<20'b00101100111001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00101100111001100110) && ({row_reg, col_reg}<20'b00101100111001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00101100111001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00101100111001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00101100111001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00101100111001101011) && ({row_reg, col_reg}<20'b00101101000100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00101101000100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00101101000100011111) && ({row_reg, col_reg}<20'b00101101000101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00101101000101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00101101000101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00101101000101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00101101000101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00101101000101010000) && ({row_reg, col_reg}<20'b00101101001000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00101101001000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00101101001000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00101101001000111000) && ({row_reg, col_reg}<20'b00101101001000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00101101001000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00101101001000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00101101001000111100) && ({row_reg, col_reg}<20'b00101101001000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00101101001000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00101101001000111111) && ({row_reg, col_reg}<20'b00101101001001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00101101001001100110) && ({row_reg, col_reg}<20'b00101101001001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00101101001001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00101101001001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00101101001001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00101101001001101011) && ({row_reg, col_reg}<20'b00101101010100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00101101010100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00101101010100011111) && ({row_reg, col_reg}<20'b00101101010101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00101101010101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00101101010101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00101101010101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00101101010101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00101101010101010000) && ({row_reg, col_reg}<20'b00101101011000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00101101011000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00101101011000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00101101011000111000) && ({row_reg, col_reg}<20'b00101101011000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00101101011000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00101101011000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00101101011000111100) && ({row_reg, col_reg}<20'b00101101011000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00101101011000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00101101011000111111) && ({row_reg, col_reg}<20'b00101101011001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00101101011001100110) && ({row_reg, col_reg}<20'b00101101011001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00101101011001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00101101011001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00101101011001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00101101011001101011) && ({row_reg, col_reg}<20'b00101101100100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00101101100100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00101101100100011111) && ({row_reg, col_reg}<20'b00101101100101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00101101100101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00101101100101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00101101100101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00101101100101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00101101100101010000) && ({row_reg, col_reg}<20'b00101101101000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00101101101000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00101101101000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00101101101000111000) && ({row_reg, col_reg}<20'b00101101101000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00101101101000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00101101101000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00101101101000111100) && ({row_reg, col_reg}<20'b00101101101000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00101101101000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00101101101000111111) && ({row_reg, col_reg}<20'b00101101101001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00101101101001100110) && ({row_reg, col_reg}<20'b00101101101001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00101101101001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00101101101001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00101101101001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00101101101001101011) && ({row_reg, col_reg}<20'b00101101110100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00101101110100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00101101110100011111) && ({row_reg, col_reg}<20'b00101101110101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00101101110101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00101101110101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00101101110101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00101101110101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00101101110101010000) && ({row_reg, col_reg}<20'b00101101111000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00101101111000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00101101111000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00101101111000111000) && ({row_reg, col_reg}<20'b00101101111000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00101101111000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00101101111000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00101101111000111100) && ({row_reg, col_reg}<20'b00101101111000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00101101111000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00101101111000111111) && ({row_reg, col_reg}<20'b00101101111001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00101101111001100110) && ({row_reg, col_reg}<20'b00101101111001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00101101111001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00101101111001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00101101111001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00101101111001101011) && ({row_reg, col_reg}<20'b00101110000100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00101110000100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00101110000100011111) && ({row_reg, col_reg}<20'b00101110000101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00101110000101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00101110000101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00101110000101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00101110000101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00101110000101010000) && ({row_reg, col_reg}<20'b00101110001000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00101110001000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00101110001000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00101110001000111000) && ({row_reg, col_reg}<20'b00101110001000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00101110001000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00101110001000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00101110001000111100) && ({row_reg, col_reg}<20'b00101110001000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00101110001000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00101110001000111111) && ({row_reg, col_reg}<20'b00101110001001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00101110001001100110) && ({row_reg, col_reg}<20'b00101110001001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00101110001001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00101110001001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00101110001001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00101110001001101011) && ({row_reg, col_reg}<20'b00101110010100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00101110010100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00101110010100011111) && ({row_reg, col_reg}<20'b00101110010101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00101110010101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00101110010101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00101110010101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00101110010101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00101110010101010000) && ({row_reg, col_reg}<20'b00101110011000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00101110011000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00101110011000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00101110011000111000) && ({row_reg, col_reg}<20'b00101110011000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00101110011000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00101110011000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00101110011000111100) && ({row_reg, col_reg}<20'b00101110011000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00101110011000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00101110011000111111) && ({row_reg, col_reg}<20'b00101110011001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00101110011001100110) && ({row_reg, col_reg}<20'b00101110011001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00101110011001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00101110011001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00101110011001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00101110011001101011) && ({row_reg, col_reg}<20'b00101110100100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00101110100100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00101110100100011111) && ({row_reg, col_reg}<20'b00101110100101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00101110100101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00101110100101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00101110100101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00101110100101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00101110100101010000) && ({row_reg, col_reg}<20'b00101110101000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00101110101000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00101110101000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00101110101000111000) && ({row_reg, col_reg}<20'b00101110101000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00101110101000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00101110101000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00101110101000111100) && ({row_reg, col_reg}<20'b00101110101000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00101110101000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00101110101000111111) && ({row_reg, col_reg}<20'b00101110101001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00101110101001100110) && ({row_reg, col_reg}<20'b00101110101001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00101110101001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00101110101001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00101110101001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00101110101001101011) && ({row_reg, col_reg}<20'b00101110110100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00101110110100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00101110110100011111) && ({row_reg, col_reg}<20'b00101110110101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00101110110101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00101110110101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00101110110101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00101110110101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00101110110101010000) && ({row_reg, col_reg}<20'b00101110111000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00101110111000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00101110111000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00101110111000111000) && ({row_reg, col_reg}<20'b00101110111000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00101110111000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00101110111000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00101110111000111100) && ({row_reg, col_reg}<20'b00101110111000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00101110111000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00101110111000111111) && ({row_reg, col_reg}<20'b00101110111001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00101110111001100110) && ({row_reg, col_reg}<20'b00101110111001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00101110111001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00101110111001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00101110111001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00101110111001101011) && ({row_reg, col_reg}<20'b00101111000100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00101111000100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00101111000100011111) && ({row_reg, col_reg}<20'b00101111000101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00101111000101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00101111000101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00101111000101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00101111000101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00101111000101010000) && ({row_reg, col_reg}<20'b00101111001000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00101111001000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00101111001000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00101111001000111000) && ({row_reg, col_reg}<20'b00101111001000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00101111001000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00101111001000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00101111001000111100) && ({row_reg, col_reg}<20'b00101111001000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00101111001000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00101111001000111111) && ({row_reg, col_reg}<20'b00101111001001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00101111001001100110) && ({row_reg, col_reg}<20'b00101111001001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00101111001001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00101111001001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00101111001001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00101111001001101011) && ({row_reg, col_reg}<20'b00101111010100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00101111010100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00101111010100011111) && ({row_reg, col_reg}<20'b00101111010101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00101111010101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00101111010101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00101111010101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00101111010101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00101111010101010000) && ({row_reg, col_reg}<20'b00101111011000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00101111011000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00101111011000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00101111011000111000) && ({row_reg, col_reg}<20'b00101111011000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00101111011000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00101111011000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00101111011000111100) && ({row_reg, col_reg}<20'b00101111011000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00101111011000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00101111011000111111) && ({row_reg, col_reg}<20'b00101111011001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00101111011001100110) && ({row_reg, col_reg}<20'b00101111011001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00101111011001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00101111011001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00101111011001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00101111011001101011) && ({row_reg, col_reg}<20'b00101111100100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00101111100100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00101111100100011111) && ({row_reg, col_reg}<20'b00101111100101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00101111100101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00101111100101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00101111100101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00101111100101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00101111100101010000) && ({row_reg, col_reg}<20'b00101111101000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00101111101000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00101111101000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00101111101000111000) && ({row_reg, col_reg}<20'b00101111101000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00101111101000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00101111101000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00101111101000111100) && ({row_reg, col_reg}<20'b00101111101000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00101111101000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00101111101000111111) && ({row_reg, col_reg}<20'b00101111101001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00101111101001100110) && ({row_reg, col_reg}<20'b00101111101001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00101111101001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00101111101001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00101111101001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00101111101001101011) && ({row_reg, col_reg}<20'b00101111110100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00101111110100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00101111110100011111) && ({row_reg, col_reg}<20'b00101111110101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00101111110101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00101111110101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00101111110101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00101111110101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00101111110101010000) && ({row_reg, col_reg}<20'b00101111111000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00101111111000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00101111111000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00101111111000111000) && ({row_reg, col_reg}<20'b00101111111000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00101111111000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00101111111000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00101111111000111100) && ({row_reg, col_reg}<20'b00101111111000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00101111111000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00101111111000111111) && ({row_reg, col_reg}<20'b00101111111001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00101111111001100110) && ({row_reg, col_reg}<20'b00101111111001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00101111111001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00101111111001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00101111111001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00101111111001101011) && ({row_reg, col_reg}<20'b00110000000100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00110000000100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00110000000100011111) && ({row_reg, col_reg}<20'b00110000000101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00110000000101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00110000000101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00110000000101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00110000000101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00110000000101010000) && ({row_reg, col_reg}<20'b00110000001000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00110000001000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00110000001000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00110000001000111000) && ({row_reg, col_reg}<20'b00110000001000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00110000001000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00110000001000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00110000001000111100) && ({row_reg, col_reg}<20'b00110000001000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00110000001000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00110000001000111111) && ({row_reg, col_reg}<20'b00110000001001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00110000001001100110) && ({row_reg, col_reg}<20'b00110000001001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00110000001001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00110000001001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00110000001001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00110000001001101011) && ({row_reg, col_reg}<20'b00110000010100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00110000010100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00110000010100011111) && ({row_reg, col_reg}<20'b00110000010101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00110000010101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00110000010101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00110000010101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00110000010101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00110000010101010000) && ({row_reg, col_reg}<20'b00110000011000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00110000011000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00110000011000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00110000011000111000) && ({row_reg, col_reg}<20'b00110000011000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00110000011000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00110000011000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00110000011000111100) && ({row_reg, col_reg}<20'b00110000011000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00110000011000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00110000011000111111) && ({row_reg, col_reg}<20'b00110000011001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00110000011001100110) && ({row_reg, col_reg}<20'b00110000011001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00110000011001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00110000011001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00110000011001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00110000011001101011) && ({row_reg, col_reg}<20'b00110000100100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00110000100100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00110000100100011111) && ({row_reg, col_reg}<20'b00110000100101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00110000100101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00110000100101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00110000100101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00110000100101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00110000100101010000) && ({row_reg, col_reg}<20'b00110000101000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00110000101000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00110000101000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00110000101000111000) && ({row_reg, col_reg}<20'b00110000101000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00110000101000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00110000101000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00110000101000111100) && ({row_reg, col_reg}<20'b00110000101000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00110000101000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00110000101000111111) && ({row_reg, col_reg}<20'b00110000101001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00110000101001100110) && ({row_reg, col_reg}<20'b00110000101001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00110000101001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00110000101001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00110000101001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00110000101001101011) && ({row_reg, col_reg}<20'b00110000110100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00110000110100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00110000110100011111) && ({row_reg, col_reg}<20'b00110000110101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00110000110101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00110000110101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00110000110101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00110000110101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00110000110101010000) && ({row_reg, col_reg}<20'b00110000111000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00110000111000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00110000111000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00110000111000111000) && ({row_reg, col_reg}<20'b00110000111000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00110000111000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00110000111000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00110000111000111100) && ({row_reg, col_reg}<20'b00110000111000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00110000111000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00110000111000111111) && ({row_reg, col_reg}<20'b00110000111001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00110000111001100110) && ({row_reg, col_reg}<20'b00110000111001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00110000111001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00110000111001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00110000111001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00110000111001101011) && ({row_reg, col_reg}<20'b00110001000100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00110001000100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00110001000100011111) && ({row_reg, col_reg}<20'b00110001000101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00110001000101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00110001000101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00110001000101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00110001000101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00110001000101010000) && ({row_reg, col_reg}<20'b00110001001000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00110001001000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00110001001000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00110001001000111000) && ({row_reg, col_reg}<20'b00110001001000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00110001001000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00110001001000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00110001001000111100) && ({row_reg, col_reg}<20'b00110001001000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00110001001000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00110001001000111111) && ({row_reg, col_reg}<20'b00110001001001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00110001001001100110) && ({row_reg, col_reg}<20'b00110001001001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00110001001001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00110001001001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00110001001001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00110001001001101011) && ({row_reg, col_reg}<20'b00110001010100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00110001010100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00110001010100011111) && ({row_reg, col_reg}<20'b00110001010101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00110001010101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00110001010101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00110001010101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00110001010101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00110001010101010000) && ({row_reg, col_reg}<20'b00110001011000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00110001011000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00110001011000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00110001011000111000) && ({row_reg, col_reg}<20'b00110001011000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00110001011000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00110001011000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00110001011000111100) && ({row_reg, col_reg}<20'b00110001011000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00110001011000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00110001011000111111) && ({row_reg, col_reg}<20'b00110001011001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00110001011001100110) && ({row_reg, col_reg}<20'b00110001011001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00110001011001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00110001011001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00110001011001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00110001011001101011) && ({row_reg, col_reg}<20'b00110001100100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00110001100100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00110001100100011111) && ({row_reg, col_reg}<20'b00110001100101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00110001100101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00110001100101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00110001100101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00110001100101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00110001100101010000) && ({row_reg, col_reg}<20'b00110001101000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00110001101000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00110001101000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00110001101000111000) && ({row_reg, col_reg}<20'b00110001101000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00110001101000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00110001101000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00110001101000111100) && ({row_reg, col_reg}<20'b00110001101000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00110001101000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00110001101000111111) && ({row_reg, col_reg}<20'b00110001101001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00110001101001100110) && ({row_reg, col_reg}<20'b00110001101001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00110001101001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00110001101001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00110001101001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00110001101001101011) && ({row_reg, col_reg}<20'b00110001110100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00110001110100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00110001110100011111) && ({row_reg, col_reg}<20'b00110001110101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00110001110101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00110001110101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00110001110101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00110001110101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00110001110101010000) && ({row_reg, col_reg}<20'b00110001111000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00110001111000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00110001111000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00110001111000111000) && ({row_reg, col_reg}<20'b00110001111000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00110001111000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00110001111000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00110001111000111100) && ({row_reg, col_reg}<20'b00110001111000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00110001111000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00110001111000111111) && ({row_reg, col_reg}<20'b00110001111001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00110001111001100110) && ({row_reg, col_reg}<20'b00110001111001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00110001111001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00110001111001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00110001111001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00110001111001101011) && ({row_reg, col_reg}<20'b00110010000100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00110010000100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00110010000100011111) && ({row_reg, col_reg}<20'b00110010000101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00110010000101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00110010000101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00110010000101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00110010000101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00110010000101010000) && ({row_reg, col_reg}<20'b00110010001000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00110010001000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00110010001000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00110010001000111000) && ({row_reg, col_reg}<20'b00110010001000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00110010001000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00110010001000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00110010001000111100) && ({row_reg, col_reg}<20'b00110010001000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00110010001000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00110010001000111111) && ({row_reg, col_reg}<20'b00110010001001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00110010001001100110) && ({row_reg, col_reg}<20'b00110010001001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00110010001001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00110010001001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00110010001001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00110010001001101011) && ({row_reg, col_reg}<20'b00110010010100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00110010010100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00110010010100011111) && ({row_reg, col_reg}<20'b00110010010101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00110010010101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00110010010101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00110010010101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00110010010101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00110010010101010000) && ({row_reg, col_reg}<20'b00110010011000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00110010011000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00110010011000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00110010011000111000) && ({row_reg, col_reg}<20'b00110010011000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00110010011000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00110010011000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00110010011000111100) && ({row_reg, col_reg}<20'b00110010011000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00110010011000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00110010011000111111) && ({row_reg, col_reg}<20'b00110010011001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00110010011001100110) && ({row_reg, col_reg}<20'b00110010011001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00110010011001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00110010011001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00110010011001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00110010011001101011) && ({row_reg, col_reg}<20'b00110010100100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00110010100100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00110010100100011111) && ({row_reg, col_reg}<20'b00110010100101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00110010100101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00110010100101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00110010100101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00110010100101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00110010100101010000) && ({row_reg, col_reg}<20'b00110010101000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00110010101000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00110010101000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00110010101000111000) && ({row_reg, col_reg}<20'b00110010101000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00110010101000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00110010101000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00110010101000111100) && ({row_reg, col_reg}<20'b00110010101000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00110010101000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00110010101000111111) && ({row_reg, col_reg}<20'b00110010101001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00110010101001100110) && ({row_reg, col_reg}<20'b00110010101001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00110010101001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00110010101001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00110010101001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00110010101001101011) && ({row_reg, col_reg}<20'b00110010110100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00110010110100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00110010110100011111) && ({row_reg, col_reg}<20'b00110010110101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00110010110101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00110010110101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00110010110101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00110010110101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00110010110101010000) && ({row_reg, col_reg}<20'b00110010111000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00110010111000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00110010111000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00110010111000111000) && ({row_reg, col_reg}<20'b00110010111000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00110010111000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00110010111000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00110010111000111100) && ({row_reg, col_reg}<20'b00110010111000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00110010111000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00110010111000111111) && ({row_reg, col_reg}<20'b00110010111001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00110010111001100110) && ({row_reg, col_reg}<20'b00110010111001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00110010111001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00110010111001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00110010111001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00110010111001101011) && ({row_reg, col_reg}<20'b00110011000100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00110011000100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00110011000100011111) && ({row_reg, col_reg}<20'b00110011000101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00110011000101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00110011000101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00110011000101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00110011000101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00110011000101010000) && ({row_reg, col_reg}<20'b00110011001000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00110011001000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00110011001000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00110011001000111000) && ({row_reg, col_reg}<20'b00110011001000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00110011001000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00110011001000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00110011001000111100) && ({row_reg, col_reg}<20'b00110011001000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00110011001000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00110011001000111111) && ({row_reg, col_reg}<20'b00110011001001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00110011001001100110) && ({row_reg, col_reg}<20'b00110011001001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00110011001001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00110011001001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00110011001001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00110011001001101011) && ({row_reg, col_reg}<20'b00110011010100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00110011010100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00110011010100011111) && ({row_reg, col_reg}<20'b00110011010101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00110011010101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00110011010101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00110011010101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00110011010101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00110011010101010000) && ({row_reg, col_reg}<20'b00110011011000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00110011011000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00110011011000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00110011011000111000) && ({row_reg, col_reg}<20'b00110011011000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00110011011000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00110011011000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00110011011000111100) && ({row_reg, col_reg}<20'b00110011011000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00110011011000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00110011011000111111) && ({row_reg, col_reg}<20'b00110011011001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00110011011001100110) && ({row_reg, col_reg}<20'b00110011011001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00110011011001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00110011011001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00110011011001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00110011011001101011) && ({row_reg, col_reg}<20'b00110011100100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00110011100100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00110011100100011111) && ({row_reg, col_reg}<20'b00110011100101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00110011100101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00110011100101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00110011100101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00110011100101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00110011100101010000) && ({row_reg, col_reg}<20'b00110011101000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00110011101000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00110011101000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00110011101000111000) && ({row_reg, col_reg}<20'b00110011101000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00110011101000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00110011101000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00110011101000111100) && ({row_reg, col_reg}<20'b00110011101000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00110011101000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00110011101000111111) && ({row_reg, col_reg}<20'b00110011101001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00110011101001100110) && ({row_reg, col_reg}<20'b00110011101001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00110011101001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00110011101001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00110011101001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00110011101001101011) && ({row_reg, col_reg}<20'b00110011110100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00110011110100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00110011110100011111) && ({row_reg, col_reg}<20'b00110011110101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00110011110101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00110011110101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00110011110101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00110011110101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00110011110101010000) && ({row_reg, col_reg}<20'b00110011111000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00110011111000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00110011111000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00110011111000111000) && ({row_reg, col_reg}<20'b00110011111000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00110011111000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00110011111000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00110011111000111100) && ({row_reg, col_reg}<20'b00110011111000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00110011111000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00110011111000111111) && ({row_reg, col_reg}<20'b00110011111001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00110011111001100110) && ({row_reg, col_reg}<20'b00110011111001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00110011111001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00110011111001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00110011111001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00110011111001101011) && ({row_reg, col_reg}<20'b00110100000100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00110100000100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00110100000100011111) && ({row_reg, col_reg}<20'b00110100000101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00110100000101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00110100000101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00110100000101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00110100000101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00110100000101010000) && ({row_reg, col_reg}<20'b00110100001000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00110100001000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00110100001000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00110100001000111000) && ({row_reg, col_reg}<20'b00110100001000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00110100001000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00110100001000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00110100001000111100) && ({row_reg, col_reg}<20'b00110100001000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00110100001000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00110100001000111111) && ({row_reg, col_reg}<20'b00110100001001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00110100001001100110) && ({row_reg, col_reg}<20'b00110100001001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00110100001001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00110100001001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00110100001001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00110100001001101011) && ({row_reg, col_reg}<20'b00110100010100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00110100010100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00110100010100011111) && ({row_reg, col_reg}<20'b00110100010101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00110100010101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00110100010101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00110100010101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00110100010101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00110100010101010000) && ({row_reg, col_reg}<20'b00110100011000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00110100011000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00110100011000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00110100011000111000) && ({row_reg, col_reg}<20'b00110100011000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00110100011000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00110100011000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00110100011000111100) && ({row_reg, col_reg}<20'b00110100011000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00110100011000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00110100011000111111) && ({row_reg, col_reg}<20'b00110100011001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00110100011001100110) && ({row_reg, col_reg}<20'b00110100011001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00110100011001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00110100011001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00110100011001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00110100011001101011) && ({row_reg, col_reg}<20'b00110100100100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00110100100100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00110100100100011111) && ({row_reg, col_reg}<20'b00110100100101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00110100100101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00110100100101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00110100100101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00110100100101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00110100100101010000) && ({row_reg, col_reg}<20'b00110100101000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00110100101000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00110100101000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00110100101000111000) && ({row_reg, col_reg}<20'b00110100101000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00110100101000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00110100101000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00110100101000111100) && ({row_reg, col_reg}<20'b00110100101000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00110100101000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00110100101000111111) && ({row_reg, col_reg}<20'b00110100101001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00110100101001100110) && ({row_reg, col_reg}<20'b00110100101001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00110100101001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00110100101001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00110100101001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00110100101001101011) && ({row_reg, col_reg}<20'b00110100110100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00110100110100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00110100110100011111) && ({row_reg, col_reg}<20'b00110100110101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00110100110101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00110100110101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00110100110101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00110100110101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00110100110101010000) && ({row_reg, col_reg}<20'b00110100111000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00110100111000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00110100111000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00110100111000111000) && ({row_reg, col_reg}<20'b00110100111000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00110100111000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00110100111000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00110100111000111100) && ({row_reg, col_reg}<20'b00110100111000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00110100111000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00110100111000111111) && ({row_reg, col_reg}<20'b00110100111001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00110100111001100110) && ({row_reg, col_reg}<20'b00110100111001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00110100111001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00110100111001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00110100111001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00110100111001101011) && ({row_reg, col_reg}<20'b00110101000100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00110101000100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00110101000100011111) && ({row_reg, col_reg}<20'b00110101000101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00110101000101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00110101000101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00110101000101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00110101000101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00110101000101010000) && ({row_reg, col_reg}<20'b00110101001000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00110101001000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00110101001000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00110101001000111000) && ({row_reg, col_reg}<20'b00110101001000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00110101001000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00110101001000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00110101001000111100) && ({row_reg, col_reg}<20'b00110101001000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00110101001000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00110101001000111111) && ({row_reg, col_reg}<20'b00110101001001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00110101001001100110) && ({row_reg, col_reg}<20'b00110101001001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00110101001001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00110101001001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00110101001001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00110101001001101011) && ({row_reg, col_reg}<20'b00110101010100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00110101010100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00110101010100011111) && ({row_reg, col_reg}<20'b00110101010101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00110101010101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00110101010101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00110101010101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00110101010101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00110101010101010000) && ({row_reg, col_reg}<20'b00110101011000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00110101011000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00110101011000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00110101011000111000) && ({row_reg, col_reg}<20'b00110101011000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00110101011000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00110101011000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00110101011000111100) && ({row_reg, col_reg}<20'b00110101011000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00110101011000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00110101011000111111) && ({row_reg, col_reg}<20'b00110101011001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00110101011001100110) && ({row_reg, col_reg}<20'b00110101011001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00110101011001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00110101011001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00110101011001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00110101011001101011) && ({row_reg, col_reg}<20'b00110101100100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00110101100100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00110101100100011111) && ({row_reg, col_reg}<20'b00110101100101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00110101100101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00110101100101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00110101100101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00110101100101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00110101100101010000) && ({row_reg, col_reg}<20'b00110101101000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00110101101000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00110101101000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00110101101000111000) && ({row_reg, col_reg}<20'b00110101101000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00110101101000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00110101101000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00110101101000111100) && ({row_reg, col_reg}<20'b00110101101000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00110101101000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00110101101000111111) && ({row_reg, col_reg}<20'b00110101101001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00110101101001100110) && ({row_reg, col_reg}<20'b00110101101001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00110101101001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00110101101001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00110101101001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00110101101001101011) && ({row_reg, col_reg}<20'b00110101110100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00110101110100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00110101110100011111) && ({row_reg, col_reg}<20'b00110101110101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00110101110101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00110101110101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00110101110101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00110101110101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00110101110101010000) && ({row_reg, col_reg}<20'b00110101111000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00110101111000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00110101111000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00110101111000111000) && ({row_reg, col_reg}<20'b00110101111000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00110101111000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00110101111000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00110101111000111100) && ({row_reg, col_reg}<20'b00110101111000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00110101111000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00110101111000111111) && ({row_reg, col_reg}<20'b00110101111001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00110101111001100110) && ({row_reg, col_reg}<20'b00110101111001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00110101111001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00110101111001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00110101111001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00110101111001101011) && ({row_reg, col_reg}<20'b00110110000100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00110110000100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00110110000100011111) && ({row_reg, col_reg}<20'b00110110000101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00110110000101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00110110000101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00110110000101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00110110000101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00110110000101010000) && ({row_reg, col_reg}<20'b00110110001000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00110110001000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00110110001000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00110110001000111000) && ({row_reg, col_reg}<20'b00110110001000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00110110001000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00110110001000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00110110001000111100) && ({row_reg, col_reg}<20'b00110110001000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00110110001000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00110110001000111111) && ({row_reg, col_reg}<20'b00110110001001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00110110001001100110) && ({row_reg, col_reg}<20'b00110110001001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00110110001001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00110110001001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00110110001001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00110110001001101011) && ({row_reg, col_reg}<20'b00110110010100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00110110010100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00110110010100011111) && ({row_reg, col_reg}<20'b00110110010101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00110110010101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00110110010101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00110110010101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00110110010101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00110110010101010000) && ({row_reg, col_reg}<20'b00110110011000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00110110011000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00110110011000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00110110011000111000) && ({row_reg, col_reg}<20'b00110110011000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00110110011000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00110110011000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00110110011000111100) && ({row_reg, col_reg}<20'b00110110011000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00110110011000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00110110011000111111) && ({row_reg, col_reg}<20'b00110110011001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00110110011001100110) && ({row_reg, col_reg}<20'b00110110011001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00110110011001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00110110011001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00110110011001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00110110011001101011) && ({row_reg, col_reg}<20'b00110110100100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00110110100100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00110110100100011111) && ({row_reg, col_reg}<20'b00110110100101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00110110100101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00110110100101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00110110100101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00110110100101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00110110100101010000) && ({row_reg, col_reg}<20'b00110110101000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00110110101000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00110110101000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00110110101000111000) && ({row_reg, col_reg}<20'b00110110101000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00110110101000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00110110101000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00110110101000111100) && ({row_reg, col_reg}<20'b00110110101000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00110110101000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00110110101000111111) && ({row_reg, col_reg}<20'b00110110101001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00110110101001100110) && ({row_reg, col_reg}<20'b00110110101001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00110110101001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00110110101001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00110110101001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00110110101001101011) && ({row_reg, col_reg}<20'b00110110110100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00110110110100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00110110110100011111) && ({row_reg, col_reg}<20'b00110110110101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00110110110101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00110110110101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00110110110101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00110110110101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00110110110101010000) && ({row_reg, col_reg}<20'b00110110111000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00110110111000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00110110111000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00110110111000111000) && ({row_reg, col_reg}<20'b00110110111000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00110110111000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00110110111000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00110110111000111100) && ({row_reg, col_reg}<20'b00110110111000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00110110111000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00110110111000111111) && ({row_reg, col_reg}<20'b00110110111001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00110110111001100110) && ({row_reg, col_reg}<20'b00110110111001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00110110111001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00110110111001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00110110111001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00110110111001101011) && ({row_reg, col_reg}<20'b00110111000100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00110111000100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00110111000100011111) && ({row_reg, col_reg}<20'b00110111000101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00110111000101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00110111000101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00110111000101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00110111000101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00110111000101010000) && ({row_reg, col_reg}<20'b00110111001000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00110111001000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00110111001000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00110111001000111000) && ({row_reg, col_reg}<20'b00110111001000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00110111001000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00110111001000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00110111001000111100) && ({row_reg, col_reg}<20'b00110111001000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00110111001000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00110111001000111111) && ({row_reg, col_reg}<20'b00110111001001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00110111001001100110) && ({row_reg, col_reg}<20'b00110111001001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00110111001001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00110111001001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00110111001001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00110111001001101011) && ({row_reg, col_reg}<20'b00110111010100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00110111010100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00110111010100011111) && ({row_reg, col_reg}<20'b00110111010101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00110111010101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00110111010101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00110111010101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00110111010101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00110111010101010000) && ({row_reg, col_reg}<20'b00110111011000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00110111011000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00110111011000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00110111011000111000) && ({row_reg, col_reg}<20'b00110111011000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00110111011000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00110111011000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00110111011000111100) && ({row_reg, col_reg}<20'b00110111011000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00110111011000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00110111011000111111) && ({row_reg, col_reg}<20'b00110111011001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00110111011001100110) && ({row_reg, col_reg}<20'b00110111011001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00110111011001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00110111011001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00110111011001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00110111011001101011) && ({row_reg, col_reg}<20'b00110111100100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00110111100100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00110111100100011111) && ({row_reg, col_reg}<20'b00110111100101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00110111100101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00110111100101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00110111100101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00110111100101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00110111100101010000) && ({row_reg, col_reg}<20'b00110111101000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00110111101000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00110111101000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00110111101000111000) && ({row_reg, col_reg}<20'b00110111101000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00110111101000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00110111101000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00110111101000111100) && ({row_reg, col_reg}<20'b00110111101000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00110111101000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00110111101000111111) && ({row_reg, col_reg}<20'b00110111101001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00110111101001100110) && ({row_reg, col_reg}<20'b00110111101001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00110111101001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00110111101001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00110111101001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00110111101001101011) && ({row_reg, col_reg}<20'b00110111110100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00110111110100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00110111110100011111) && ({row_reg, col_reg}<20'b00110111110101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00110111110101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00110111110101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00110111110101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00110111110101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00110111110101010000) && ({row_reg, col_reg}<20'b00110111111000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00110111111000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00110111111000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00110111111000111000) && ({row_reg, col_reg}<20'b00110111111000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00110111111000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00110111111000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00110111111000111100) && ({row_reg, col_reg}<20'b00110111111000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00110111111000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00110111111000111111) && ({row_reg, col_reg}<20'b00110111111001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00110111111001100110) && ({row_reg, col_reg}<20'b00110111111001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00110111111001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00110111111001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00110111111001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00110111111001101011) && ({row_reg, col_reg}<20'b00111000000100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00111000000100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00111000000100011111) && ({row_reg, col_reg}<20'b00111000000101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00111000000101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00111000000101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00111000000101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00111000000101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00111000000101010000) && ({row_reg, col_reg}<20'b00111000001000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00111000001000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00111000001000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00111000001000111000) && ({row_reg, col_reg}<20'b00111000001000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00111000001000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00111000001000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00111000001000111100) && ({row_reg, col_reg}<20'b00111000001000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00111000001000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00111000001000111111) && ({row_reg, col_reg}<20'b00111000001001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00111000001001100110) && ({row_reg, col_reg}<20'b00111000001001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00111000001001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00111000001001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00111000001001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00111000001001101011) && ({row_reg, col_reg}<20'b00111000010100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00111000010100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00111000010100011111) && ({row_reg, col_reg}<20'b00111000010101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00111000010101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00111000010101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00111000010101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00111000010101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00111000010101010000) && ({row_reg, col_reg}<20'b00111000011000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00111000011000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00111000011000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00111000011000111000) && ({row_reg, col_reg}<20'b00111000011000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00111000011000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00111000011000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00111000011000111100) && ({row_reg, col_reg}<20'b00111000011000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00111000011000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00111000011000111111) && ({row_reg, col_reg}<20'b00111000011001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00111000011001100110) && ({row_reg, col_reg}<20'b00111000011001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00111000011001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00111000011001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00111000011001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00111000011001101011) && ({row_reg, col_reg}<20'b00111000100100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00111000100100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00111000100100011111) && ({row_reg, col_reg}<20'b00111000100101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00111000100101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00111000100101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00111000100101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00111000100101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00111000100101010000) && ({row_reg, col_reg}<20'b00111000101000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00111000101000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00111000101000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00111000101000111000) && ({row_reg, col_reg}<20'b00111000101000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00111000101000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00111000101000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00111000101000111100) && ({row_reg, col_reg}<20'b00111000101000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00111000101000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00111000101000111111) && ({row_reg, col_reg}<20'b00111000101001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00111000101001100110) && ({row_reg, col_reg}<20'b00111000101001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00111000101001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00111000101001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00111000101001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00111000101001101011) && ({row_reg, col_reg}<20'b00111000110100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00111000110100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00111000110100011111) && ({row_reg, col_reg}<20'b00111000110101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00111000110101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00111000110101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00111000110101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00111000110101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00111000110101010000) && ({row_reg, col_reg}<20'b00111000111000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00111000111000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00111000111000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00111000111000111000) && ({row_reg, col_reg}<20'b00111000111000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00111000111000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00111000111000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00111000111000111100) && ({row_reg, col_reg}<20'b00111000111000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00111000111000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00111000111000111111) && ({row_reg, col_reg}<20'b00111000111001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00111000111001100110) && ({row_reg, col_reg}<20'b00111000111001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00111000111001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00111000111001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00111000111001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00111000111001101011) && ({row_reg, col_reg}<20'b00111001000100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00111001000100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00111001000100011111) && ({row_reg, col_reg}<20'b00111001000101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00111001000101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00111001000101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00111001000101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00111001000101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00111001000101010000) && ({row_reg, col_reg}<20'b00111001001000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00111001001000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00111001001000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00111001001000111000) && ({row_reg, col_reg}<20'b00111001001000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00111001001000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00111001001000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00111001001000111100) && ({row_reg, col_reg}<20'b00111001001000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00111001001000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00111001001000111111) && ({row_reg, col_reg}<20'b00111001001001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00111001001001100110) && ({row_reg, col_reg}<20'b00111001001001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00111001001001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00111001001001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00111001001001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00111001001001101011) && ({row_reg, col_reg}<20'b00111001010100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00111001010100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00111001010100011111) && ({row_reg, col_reg}<20'b00111001010101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00111001010101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00111001010101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00111001010101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00111001010101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00111001010101010000) && ({row_reg, col_reg}<20'b00111001011000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00111001011000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00111001011000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00111001011000111000) && ({row_reg, col_reg}<20'b00111001011000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00111001011000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00111001011000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00111001011000111100) && ({row_reg, col_reg}<20'b00111001011000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00111001011000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00111001011000111111) && ({row_reg, col_reg}<20'b00111001011001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00111001011001100110) && ({row_reg, col_reg}<20'b00111001011001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00111001011001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00111001011001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00111001011001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00111001011001101011) && ({row_reg, col_reg}<20'b00111001100100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00111001100100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00111001100100011111) && ({row_reg, col_reg}<20'b00111001100101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00111001100101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00111001100101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00111001100101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00111001100101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00111001100101010000) && ({row_reg, col_reg}<20'b00111001101000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00111001101000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00111001101000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00111001101000111000) && ({row_reg, col_reg}<20'b00111001101000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00111001101000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00111001101000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00111001101000111100) && ({row_reg, col_reg}<20'b00111001101000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00111001101000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00111001101000111111) && ({row_reg, col_reg}<20'b00111001101001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00111001101001100110) && ({row_reg, col_reg}<20'b00111001101001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00111001101001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00111001101001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00111001101001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00111001101001101011) && ({row_reg, col_reg}<20'b00111001110100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00111001110100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00111001110100011111) && ({row_reg, col_reg}<20'b00111001110101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00111001110101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00111001110101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00111001110101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00111001110101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00111001110101010000) && ({row_reg, col_reg}<20'b00111001111000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00111001111000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00111001111000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00111001111000111000) && ({row_reg, col_reg}<20'b00111001111000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00111001111000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00111001111000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00111001111000111100) && ({row_reg, col_reg}<20'b00111001111000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00111001111000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00111001111000111111) && ({row_reg, col_reg}<20'b00111001111001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00111001111001100110) && ({row_reg, col_reg}<20'b00111001111001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00111001111001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00111001111001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00111001111001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00111001111001101011) && ({row_reg, col_reg}<20'b00111010000100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00111010000100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00111010000100011111) && ({row_reg, col_reg}<20'b00111010000101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00111010000101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00111010000101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00111010000101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00111010000101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00111010000101010000) && ({row_reg, col_reg}<20'b00111010001000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00111010001000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00111010001000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00111010001000111000) && ({row_reg, col_reg}<20'b00111010001000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00111010001000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00111010001000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00111010001000111100) && ({row_reg, col_reg}<20'b00111010001000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00111010001000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00111010001000111111) && ({row_reg, col_reg}<20'b00111010001001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00111010001001100110) && ({row_reg, col_reg}<20'b00111010001001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00111010001001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00111010001001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00111010001001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00111010001001101011) && ({row_reg, col_reg}<20'b00111010010100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00111010010100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00111010010100011111) && ({row_reg, col_reg}<20'b00111010010101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00111010010101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00111010010101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00111010010101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00111010010101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00111010010101010000) && ({row_reg, col_reg}<20'b00111010011000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00111010011000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00111010011000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00111010011000111000) && ({row_reg, col_reg}<20'b00111010011000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00111010011000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00111010011000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00111010011000111100) && ({row_reg, col_reg}<20'b00111010011000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00111010011000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00111010011000111111) && ({row_reg, col_reg}<20'b00111010011001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00111010011001100110) && ({row_reg, col_reg}<20'b00111010011001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00111010011001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00111010011001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00111010011001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00111010011001101011) && ({row_reg, col_reg}<20'b00111010100100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00111010100100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00111010100100011111) && ({row_reg, col_reg}<20'b00111010100101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00111010100101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00111010100101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00111010100101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00111010100101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00111010100101010000) && ({row_reg, col_reg}<20'b00111010101000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00111010101000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00111010101000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00111010101000111000) && ({row_reg, col_reg}<20'b00111010101000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00111010101000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00111010101000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00111010101000111100) && ({row_reg, col_reg}<20'b00111010101000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00111010101000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00111010101000111111) && ({row_reg, col_reg}<20'b00111010101001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00111010101001100110) && ({row_reg, col_reg}<20'b00111010101001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00111010101001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00111010101001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00111010101001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00111010101001101011) && ({row_reg, col_reg}<20'b00111010110100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00111010110100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00111010110100011111) && ({row_reg, col_reg}<20'b00111010110101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00111010110101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00111010110101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00111010110101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00111010110101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00111010110101010000) && ({row_reg, col_reg}<20'b00111010111000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00111010111000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00111010111000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00111010111000111000) && ({row_reg, col_reg}<20'b00111010111000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00111010111000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00111010111000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00111010111000111100) && ({row_reg, col_reg}<20'b00111010111000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00111010111000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00111010111000111111) && ({row_reg, col_reg}<20'b00111010111001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00111010111001100110) && ({row_reg, col_reg}<20'b00111010111001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00111010111001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00111010111001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00111010111001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00111010111001101011) && ({row_reg, col_reg}<20'b00111011000100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00111011000100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00111011000100011111) && ({row_reg, col_reg}<20'b00111011000101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00111011000101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00111011000101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00111011000101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00111011000101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00111011000101010000) && ({row_reg, col_reg}<20'b00111011001000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00111011001000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00111011001000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00111011001000111000) && ({row_reg, col_reg}<20'b00111011001000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00111011001000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00111011001000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00111011001000111100) && ({row_reg, col_reg}<20'b00111011001000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00111011001000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00111011001000111111) && ({row_reg, col_reg}<20'b00111011001001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00111011001001100110) && ({row_reg, col_reg}<20'b00111011001001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00111011001001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00111011001001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00111011001001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00111011001001101011) && ({row_reg, col_reg}<20'b00111011010100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00111011010100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00111011010100011111) && ({row_reg, col_reg}<20'b00111011010101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00111011010101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00111011010101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00111011010101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00111011010101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00111011010101010000) && ({row_reg, col_reg}<20'b00111011011000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00111011011000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00111011011000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00111011011000111000) && ({row_reg, col_reg}<20'b00111011011000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00111011011000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00111011011000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00111011011000111100) && ({row_reg, col_reg}<20'b00111011011000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00111011011000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00111011011000111111) && ({row_reg, col_reg}<20'b00111011011001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00111011011001100110) && ({row_reg, col_reg}<20'b00111011011001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00111011011001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00111011011001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00111011011001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00111011011001101011) && ({row_reg, col_reg}<20'b00111011100100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00111011100100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00111011100100011111) && ({row_reg, col_reg}<20'b00111011100101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00111011100101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00111011100101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00111011100101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00111011100101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00111011100101010000) && ({row_reg, col_reg}<20'b00111011101000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00111011101000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00111011101000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00111011101000111000) && ({row_reg, col_reg}<20'b00111011101000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00111011101000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00111011101000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00111011101000111100) && ({row_reg, col_reg}<20'b00111011101000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00111011101000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00111011101000111111) && ({row_reg, col_reg}<20'b00111011101001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00111011101001100110) && ({row_reg, col_reg}<20'b00111011101001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00111011101001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00111011101001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00111011101001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00111011101001101011) && ({row_reg, col_reg}<20'b00111011110100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00111011110100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00111011110100011111) && ({row_reg, col_reg}<20'b00111011110101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00111011110101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00111011110101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00111011110101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00111011110101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00111011110101010000) && ({row_reg, col_reg}<20'b00111011111000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00111011111000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00111011111000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00111011111000111000) && ({row_reg, col_reg}<20'b00111011111000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00111011111000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00111011111000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00111011111000111100) && ({row_reg, col_reg}<20'b00111011111000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00111011111000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00111011111000111111) && ({row_reg, col_reg}<20'b00111011111001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00111011111001100110) && ({row_reg, col_reg}<20'b00111011111001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00111011111001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00111011111001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00111011111001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00111011111001101011) && ({row_reg, col_reg}<20'b00111100000100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00111100000100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00111100000100011111) && ({row_reg, col_reg}<20'b00111100000101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00111100000101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00111100000101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00111100000101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00111100000101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00111100000101010000) && ({row_reg, col_reg}<20'b00111100001000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00111100001000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00111100001000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00111100001000111000) && ({row_reg, col_reg}<20'b00111100001000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00111100001000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00111100001000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00111100001000111100) && ({row_reg, col_reg}<20'b00111100001000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00111100001000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00111100001000111111) && ({row_reg, col_reg}<20'b00111100001001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00111100001001100110) && ({row_reg, col_reg}<20'b00111100001001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00111100001001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00111100001001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00111100001001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00111100001001101011) && ({row_reg, col_reg}<20'b00111100010100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00111100010100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00111100010100011111) && ({row_reg, col_reg}<20'b00111100010101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00111100010101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00111100010101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00111100010101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00111100010101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00111100010101010000) && ({row_reg, col_reg}<20'b00111100011000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00111100011000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00111100011000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00111100011000111000) && ({row_reg, col_reg}<20'b00111100011000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00111100011000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00111100011000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00111100011000111100) && ({row_reg, col_reg}<20'b00111100011000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00111100011000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00111100011000111111) && ({row_reg, col_reg}<20'b00111100011001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00111100011001100110) && ({row_reg, col_reg}<20'b00111100011001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00111100011001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00111100011001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00111100011001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00111100011001101011) && ({row_reg, col_reg}<20'b00111100100100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00111100100100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00111100100100011111) && ({row_reg, col_reg}<20'b00111100100101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00111100100101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00111100100101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00111100100101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00111100100101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00111100100101010000) && ({row_reg, col_reg}<20'b00111100101000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00111100101000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00111100101000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00111100101000111000) && ({row_reg, col_reg}<20'b00111100101000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00111100101000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00111100101000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00111100101000111100) && ({row_reg, col_reg}<20'b00111100101000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00111100101000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00111100101000111111) && ({row_reg, col_reg}<20'b00111100101001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00111100101001100110) && ({row_reg, col_reg}<20'b00111100101001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00111100101001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00111100101001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00111100101001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00111100101001101011) && ({row_reg, col_reg}<20'b00111100110100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00111100110100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00111100110100011111) && ({row_reg, col_reg}<20'b00111100110101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00111100110101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00111100110101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00111100110101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00111100110101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00111100110101010000) && ({row_reg, col_reg}<20'b00111100111000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00111100111000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00111100111000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00111100111000111000) && ({row_reg, col_reg}<20'b00111100111000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00111100111000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00111100111000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00111100111000111100) && ({row_reg, col_reg}<20'b00111100111000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00111100111000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00111100111000111111) && ({row_reg, col_reg}<20'b00111100111001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00111100111001100110) && ({row_reg, col_reg}<20'b00111100111001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00111100111001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00111100111001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00111100111001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00111100111001101011) && ({row_reg, col_reg}<20'b00111101000100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00111101000100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00111101000100011111) && ({row_reg, col_reg}<20'b00111101000101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00111101000101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00111101000101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00111101000101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00111101000101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00111101000101010000) && ({row_reg, col_reg}<20'b00111101001000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00111101001000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00111101001000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00111101001000111000) && ({row_reg, col_reg}<20'b00111101001000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00111101001000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00111101001000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00111101001000111100) && ({row_reg, col_reg}<20'b00111101001000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00111101001000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00111101001000111111) && ({row_reg, col_reg}<20'b00111101001001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00111101001001100110) && ({row_reg, col_reg}<20'b00111101001001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00111101001001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00111101001001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00111101001001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00111101001001101011) && ({row_reg, col_reg}<20'b00111101010100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00111101010100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00111101010100011111) && ({row_reg, col_reg}<20'b00111101010101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00111101010101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00111101010101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00111101010101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00111101010101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00111101010101010000) && ({row_reg, col_reg}<20'b00111101011000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00111101011000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00111101011000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00111101011000111000) && ({row_reg, col_reg}<20'b00111101011000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00111101011000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00111101011000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00111101011000111100) && ({row_reg, col_reg}<20'b00111101011000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00111101011000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00111101011000111111) && ({row_reg, col_reg}<20'b00111101011001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00111101011001100110) && ({row_reg, col_reg}<20'b00111101011001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00111101011001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00111101011001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00111101011001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00111101011001101011) && ({row_reg, col_reg}<20'b00111101100100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00111101100100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00111101100100011111) && ({row_reg, col_reg}<20'b00111101100101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00111101100101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00111101100101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00111101100101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00111101100101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00111101100101010000) && ({row_reg, col_reg}<20'b00111101101000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00111101101000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00111101101000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00111101101000111000) && ({row_reg, col_reg}<20'b00111101101000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00111101101000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00111101101000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00111101101000111100) && ({row_reg, col_reg}<20'b00111101101000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00111101101000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00111101101000111111) && ({row_reg, col_reg}<20'b00111101101001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00111101101001100110) && ({row_reg, col_reg}<20'b00111101101001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00111101101001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00111101101001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00111101101001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00111101101001101011) && ({row_reg, col_reg}<20'b00111101110100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00111101110100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00111101110100011111) && ({row_reg, col_reg}<20'b00111101110101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00111101110101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00111101110101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00111101110101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00111101110101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00111101110101010000) && ({row_reg, col_reg}<20'b00111101111000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00111101111000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00111101111000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00111101111000111000) && ({row_reg, col_reg}<20'b00111101111000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00111101111000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00111101111000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00111101111000111100) && ({row_reg, col_reg}<20'b00111101111000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00111101111000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00111101111000111111) && ({row_reg, col_reg}<20'b00111101111001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00111101111001100110) && ({row_reg, col_reg}<20'b00111101111001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00111101111001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00111101111001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00111101111001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00111101111001101011) && ({row_reg, col_reg}<20'b00111110000100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00111110000100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00111110000100011111) && ({row_reg, col_reg}<20'b00111110000101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00111110000101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00111110000101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00111110000101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00111110000101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00111110000101010000) && ({row_reg, col_reg}<20'b00111110001000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00111110001000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00111110001000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00111110001000111000) && ({row_reg, col_reg}<20'b00111110001000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00111110001000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00111110001000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00111110001000111100) && ({row_reg, col_reg}<20'b00111110001000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00111110001000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00111110001000111111) && ({row_reg, col_reg}<20'b00111110001001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00111110001001100110) && ({row_reg, col_reg}<20'b00111110001001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00111110001001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00111110001001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00111110001001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00111110001001101011) && ({row_reg, col_reg}<20'b00111110010100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00111110010100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00111110010100011111) && ({row_reg, col_reg}<20'b00111110010101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00111110010101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00111110010101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00111110010101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00111110010101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00111110010101010000) && ({row_reg, col_reg}<20'b00111110011000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00111110011000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00111110011000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00111110011000111000) && ({row_reg, col_reg}<20'b00111110011000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00111110011000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00111110011000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00111110011000111100) && ({row_reg, col_reg}<20'b00111110011000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00111110011000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00111110011000111111) && ({row_reg, col_reg}<20'b00111110011001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00111110011001100110) && ({row_reg, col_reg}<20'b00111110011001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00111110011001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00111110011001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00111110011001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00111110011001101011) && ({row_reg, col_reg}<20'b00111110100100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00111110100100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00111110100100011111) && ({row_reg, col_reg}<20'b00111110100101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00111110100101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00111110100101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00111110100101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00111110100101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00111110100101010000) && ({row_reg, col_reg}<20'b00111110101000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00111110101000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00111110101000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00111110101000111000) && ({row_reg, col_reg}<20'b00111110101000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00111110101000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00111110101000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00111110101000111100) && ({row_reg, col_reg}<20'b00111110101000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00111110101000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00111110101000111111) && ({row_reg, col_reg}<20'b00111110101001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00111110101001100110) && ({row_reg, col_reg}<20'b00111110101001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00111110101001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00111110101001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00111110101001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00111110101001101011) && ({row_reg, col_reg}<20'b00111110110100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00111110110100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00111110110100011111) && ({row_reg, col_reg}<20'b00111110110101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00111110110101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00111110110101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00111110110101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00111110110101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00111110110101010000) && ({row_reg, col_reg}<20'b00111110111000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00111110111000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00111110111000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00111110111000111000) && ({row_reg, col_reg}<20'b00111110111000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00111110111000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00111110111000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00111110111000111100) && ({row_reg, col_reg}<20'b00111110111000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00111110111000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00111110111000111111) && ({row_reg, col_reg}<20'b00111110111001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00111110111001100110) && ({row_reg, col_reg}<20'b00111110111001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00111110111001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00111110111001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00111110111001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00111110111001101011) && ({row_reg, col_reg}<20'b00111111000100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00111111000100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00111111000100011111) && ({row_reg, col_reg}<20'b00111111000101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00111111000101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00111111000101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00111111000101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00111111000101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00111111000101010000) && ({row_reg, col_reg}<20'b00111111001000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00111111001000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00111111001000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00111111001000111000) && ({row_reg, col_reg}<20'b00111111001000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00111111001000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00111111001000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00111111001000111100) && ({row_reg, col_reg}<20'b00111111001000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00111111001000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00111111001000111111) && ({row_reg, col_reg}<20'b00111111001001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00111111001001100110) && ({row_reg, col_reg}<20'b00111111001001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00111111001001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00111111001001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00111111001001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00111111001001101011) && ({row_reg, col_reg}<20'b00111111010100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00111111010100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00111111010100011111) && ({row_reg, col_reg}<20'b00111111010101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00111111010101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00111111010101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00111111010101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00111111010101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00111111010101010000) && ({row_reg, col_reg}<20'b00111111011000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00111111011000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00111111011000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00111111011000111000) && ({row_reg, col_reg}<20'b00111111011000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00111111011000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00111111011000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00111111011000111100) && ({row_reg, col_reg}<20'b00111111011000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00111111011000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00111111011000111111) && ({row_reg, col_reg}<20'b00111111011001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00111111011001100110) && ({row_reg, col_reg}<20'b00111111011001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00111111011001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00111111011001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00111111011001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00111111011001101011) && ({row_reg, col_reg}<20'b00111111100100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00111111100100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00111111100100011111) && ({row_reg, col_reg}<20'b00111111100101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00111111100101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00111111100101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00111111100101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00111111100101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00111111100101010000) && ({row_reg, col_reg}<20'b00111111101000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00111111101000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00111111101000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00111111101000111000) && ({row_reg, col_reg}<20'b00111111101000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00111111101000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00111111101000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00111111101000111100) && ({row_reg, col_reg}<20'b00111111101000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00111111101000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00111111101000111111) && ({row_reg, col_reg}<20'b00111111101001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00111111101001100110) && ({row_reg, col_reg}<20'b00111111101001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00111111101001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00111111101001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00111111101001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00111111101001101011) && ({row_reg, col_reg}<20'b00111111110100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00111111110100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b00111111110100011111) && ({row_reg, col_reg}<20'b00111111110101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00111111110101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00111111110101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00111111110101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00111111110101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00111111110101010000) && ({row_reg, col_reg}<20'b00111111111000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00111111111000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b00111111111000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b00111111111000111000) && ({row_reg, col_reg}<20'b00111111111000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00111111111000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00111111111000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00111111111000111100) && ({row_reg, col_reg}<20'b00111111111000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b00111111111000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b00111111111000111111) && ({row_reg, col_reg}<20'b00111111111001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b00111111111001100110) && ({row_reg, col_reg}<20'b00111111111001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b00111111111001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b00111111111001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b00111111111001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b00111111111001101011) && ({row_reg, col_reg}<20'b01000000000100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01000000000100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01000000000100011111) && ({row_reg, col_reg}<20'b01000000000101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01000000000101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01000000000101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01000000000101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01000000000101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01000000000101010000) && ({row_reg, col_reg}<20'b01000000001000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01000000001000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01000000001000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01000000001000111000) && ({row_reg, col_reg}<20'b01000000001000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01000000001000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01000000001000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01000000001000111100) && ({row_reg, col_reg}<20'b01000000001000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01000000001000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01000000001000111111) && ({row_reg, col_reg}<20'b01000000001001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01000000001001100110) && ({row_reg, col_reg}<20'b01000000001001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01000000001001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01000000001001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01000000001001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01000000001001101011) && ({row_reg, col_reg}<20'b01000000010100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01000000010100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01000000010100011111) && ({row_reg, col_reg}<20'b01000000010101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01000000010101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01000000010101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01000000010101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01000000010101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01000000010101010000) && ({row_reg, col_reg}<20'b01000000011000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01000000011000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01000000011000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01000000011000111000) && ({row_reg, col_reg}<20'b01000000011000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01000000011000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01000000011000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01000000011000111100) && ({row_reg, col_reg}<20'b01000000011000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01000000011000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01000000011000111111) && ({row_reg, col_reg}<20'b01000000011001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01000000011001100110) && ({row_reg, col_reg}<20'b01000000011001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01000000011001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01000000011001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01000000011001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01000000011001101011) && ({row_reg, col_reg}<20'b01000000100100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01000000100100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01000000100100011111) && ({row_reg, col_reg}<20'b01000000100101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01000000100101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01000000100101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01000000100101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01000000100101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01000000100101010000) && ({row_reg, col_reg}<20'b01000000101000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01000000101000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01000000101000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01000000101000111000) && ({row_reg, col_reg}<20'b01000000101000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01000000101000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01000000101000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01000000101000111100) && ({row_reg, col_reg}<20'b01000000101000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01000000101000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01000000101000111111) && ({row_reg, col_reg}<20'b01000000101001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01000000101001100110) && ({row_reg, col_reg}<20'b01000000101001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01000000101001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01000000101001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01000000101001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01000000101001101011) && ({row_reg, col_reg}<20'b01000000110100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01000000110100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01000000110100011111) && ({row_reg, col_reg}<20'b01000000110101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01000000110101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01000000110101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01000000110101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01000000110101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01000000110101010000) && ({row_reg, col_reg}<20'b01000000111000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01000000111000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01000000111000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01000000111000111000) && ({row_reg, col_reg}<20'b01000000111000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01000000111000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01000000111000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01000000111000111100) && ({row_reg, col_reg}<20'b01000000111000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01000000111000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01000000111000111111) && ({row_reg, col_reg}<20'b01000000111001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01000000111001100110) && ({row_reg, col_reg}<20'b01000000111001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01000000111001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01000000111001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01000000111001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01000000111001101011) && ({row_reg, col_reg}<20'b01000001000100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01000001000100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01000001000100011111) && ({row_reg, col_reg}<20'b01000001000101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01000001000101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01000001000101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01000001000101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01000001000101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01000001000101010000) && ({row_reg, col_reg}<20'b01000001001000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01000001001000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01000001001000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01000001001000111000) && ({row_reg, col_reg}<20'b01000001001000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01000001001000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01000001001000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01000001001000111100) && ({row_reg, col_reg}<20'b01000001001000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01000001001000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01000001001000111111) && ({row_reg, col_reg}<20'b01000001001001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01000001001001100110) && ({row_reg, col_reg}<20'b01000001001001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01000001001001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01000001001001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01000001001001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01000001001001101011) && ({row_reg, col_reg}<20'b01000001010100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01000001010100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01000001010100011111) && ({row_reg, col_reg}<20'b01000001010101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01000001010101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01000001010101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01000001010101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01000001010101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01000001010101010000) && ({row_reg, col_reg}<20'b01000001011000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01000001011000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01000001011000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01000001011000111000) && ({row_reg, col_reg}<20'b01000001011000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01000001011000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01000001011000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01000001011000111100) && ({row_reg, col_reg}<20'b01000001011000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01000001011000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01000001011000111111) && ({row_reg, col_reg}<20'b01000001011001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01000001011001100110) && ({row_reg, col_reg}<20'b01000001011001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01000001011001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01000001011001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01000001011001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01000001011001101011) && ({row_reg, col_reg}<20'b01000001100100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01000001100100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01000001100100011111) && ({row_reg, col_reg}<20'b01000001100101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01000001100101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01000001100101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01000001100101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01000001100101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01000001100101010000) && ({row_reg, col_reg}<20'b01000001101000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01000001101000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01000001101000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01000001101000111000) && ({row_reg, col_reg}<20'b01000001101000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01000001101000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01000001101000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01000001101000111100) && ({row_reg, col_reg}<20'b01000001101000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01000001101000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01000001101000111111) && ({row_reg, col_reg}<20'b01000001101001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01000001101001100110) && ({row_reg, col_reg}<20'b01000001101001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01000001101001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01000001101001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01000001101001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01000001101001101011) && ({row_reg, col_reg}<20'b01000001110100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01000001110100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01000001110100011111) && ({row_reg, col_reg}<20'b01000001110101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01000001110101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01000001110101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01000001110101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01000001110101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01000001110101010000) && ({row_reg, col_reg}<20'b01000001111000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01000001111000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01000001111000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01000001111000111000) && ({row_reg, col_reg}<20'b01000001111000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01000001111000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01000001111000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01000001111000111100) && ({row_reg, col_reg}<20'b01000001111000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01000001111000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01000001111000111111) && ({row_reg, col_reg}<20'b01000001111001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01000001111001100110) && ({row_reg, col_reg}<20'b01000001111001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01000001111001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01000001111001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01000001111001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01000001111001101011) && ({row_reg, col_reg}<20'b01000010000100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01000010000100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01000010000100011111) && ({row_reg, col_reg}<20'b01000010000101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01000010000101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01000010000101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01000010000101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01000010000101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01000010000101010000) && ({row_reg, col_reg}<20'b01000010001000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01000010001000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01000010001000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01000010001000111000) && ({row_reg, col_reg}<20'b01000010001000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01000010001000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01000010001000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01000010001000111100) && ({row_reg, col_reg}<20'b01000010001000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01000010001000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01000010001000111111) && ({row_reg, col_reg}<20'b01000010001001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01000010001001100110) && ({row_reg, col_reg}<20'b01000010001001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01000010001001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01000010001001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01000010001001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01000010001001101011) && ({row_reg, col_reg}<20'b01000010010100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01000010010100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01000010010100011111) && ({row_reg, col_reg}<20'b01000010010101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01000010010101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01000010010101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01000010010101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01000010010101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01000010010101010000) && ({row_reg, col_reg}<20'b01000010011000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01000010011000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01000010011000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01000010011000111000) && ({row_reg, col_reg}<20'b01000010011000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01000010011000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01000010011000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01000010011000111100) && ({row_reg, col_reg}<20'b01000010011000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01000010011000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01000010011000111111) && ({row_reg, col_reg}<20'b01000010011001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01000010011001100110) && ({row_reg, col_reg}<20'b01000010011001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01000010011001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01000010011001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01000010011001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01000010011001101011) && ({row_reg, col_reg}<20'b01000010100100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01000010100100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01000010100100011111) && ({row_reg, col_reg}<20'b01000010100101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01000010100101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01000010100101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01000010100101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01000010100101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01000010100101010000) && ({row_reg, col_reg}<20'b01000010101000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01000010101000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01000010101000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01000010101000111000) && ({row_reg, col_reg}<20'b01000010101000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01000010101000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01000010101000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01000010101000111100) && ({row_reg, col_reg}<20'b01000010101000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01000010101000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01000010101000111111) && ({row_reg, col_reg}<20'b01000010101001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01000010101001100110) && ({row_reg, col_reg}<20'b01000010101001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01000010101001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01000010101001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01000010101001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01000010101001101011) && ({row_reg, col_reg}<20'b01000010110100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01000010110100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01000010110100011111) && ({row_reg, col_reg}<20'b01000010110101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01000010110101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01000010110101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01000010110101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01000010110101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01000010110101010000) && ({row_reg, col_reg}<20'b01000010111000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01000010111000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01000010111000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01000010111000111000) && ({row_reg, col_reg}<20'b01000010111000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01000010111000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01000010111000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01000010111000111100) && ({row_reg, col_reg}<20'b01000010111000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01000010111000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01000010111000111111) && ({row_reg, col_reg}<20'b01000010111001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01000010111001100110) && ({row_reg, col_reg}<20'b01000010111001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01000010111001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01000010111001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01000010111001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01000010111001101011) && ({row_reg, col_reg}<20'b01000011000100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01000011000100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01000011000100011111) && ({row_reg, col_reg}<20'b01000011000101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01000011000101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01000011000101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01000011000101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01000011000101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01000011000101010000) && ({row_reg, col_reg}<20'b01000011001000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01000011001000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01000011001000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01000011001000111000) && ({row_reg, col_reg}<20'b01000011001000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01000011001000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01000011001000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01000011001000111100) && ({row_reg, col_reg}<20'b01000011001000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01000011001000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01000011001000111111) && ({row_reg, col_reg}<20'b01000011001001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01000011001001100110) && ({row_reg, col_reg}<20'b01000011001001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01000011001001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01000011001001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01000011001001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01000011001001101011) && ({row_reg, col_reg}<20'b01000011010100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01000011010100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01000011010100011111) && ({row_reg, col_reg}<20'b01000011010101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01000011010101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01000011010101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01000011010101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01000011010101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01000011010101010000) && ({row_reg, col_reg}<20'b01000011011000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01000011011000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01000011011000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01000011011000111000) && ({row_reg, col_reg}<20'b01000011011000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01000011011000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01000011011000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01000011011000111100) && ({row_reg, col_reg}<20'b01000011011000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01000011011000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01000011011000111111) && ({row_reg, col_reg}<20'b01000011011001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01000011011001100110) && ({row_reg, col_reg}<20'b01000011011001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01000011011001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01000011011001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01000011011001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01000011011001101011) && ({row_reg, col_reg}<20'b01000011100100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01000011100100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01000011100100011111) && ({row_reg, col_reg}<20'b01000011100101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01000011100101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01000011100101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01000011100101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01000011100101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01000011100101010000) && ({row_reg, col_reg}<20'b01000011101000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01000011101000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01000011101000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01000011101000111000) && ({row_reg, col_reg}<20'b01000011101000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01000011101000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01000011101000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01000011101000111100) && ({row_reg, col_reg}<20'b01000011101000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01000011101000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01000011101000111111) && ({row_reg, col_reg}<20'b01000011101001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01000011101001100110) && ({row_reg, col_reg}<20'b01000011101001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01000011101001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01000011101001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01000011101001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01000011101001101011) && ({row_reg, col_reg}<20'b01000011110100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01000011110100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01000011110100011111) && ({row_reg, col_reg}<20'b01000011110101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01000011110101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01000011110101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01000011110101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01000011110101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01000011110101010000) && ({row_reg, col_reg}<20'b01000011111000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01000011111000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01000011111000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01000011111000111000) && ({row_reg, col_reg}<20'b01000011111000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01000011111000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01000011111000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01000011111000111100) && ({row_reg, col_reg}<20'b01000011111000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01000011111000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01000011111000111111) && ({row_reg, col_reg}<20'b01000011111001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01000011111001100110) && ({row_reg, col_reg}<20'b01000011111001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01000011111001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01000011111001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01000011111001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01000011111001101011) && ({row_reg, col_reg}<20'b01000100000100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01000100000100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01000100000100011111) && ({row_reg, col_reg}<20'b01000100000101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01000100000101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01000100000101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01000100000101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01000100000101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01000100000101010000) && ({row_reg, col_reg}<20'b01000100001000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01000100001000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01000100001000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01000100001000111000) && ({row_reg, col_reg}<20'b01000100001000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01000100001000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01000100001000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01000100001000111100) && ({row_reg, col_reg}<20'b01000100001000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01000100001000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01000100001000111111) && ({row_reg, col_reg}<20'b01000100001001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01000100001001100110) && ({row_reg, col_reg}<20'b01000100001001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01000100001001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01000100001001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01000100001001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01000100001001101011) && ({row_reg, col_reg}<20'b01000100010100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01000100010100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01000100010100011111) && ({row_reg, col_reg}<20'b01000100010101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01000100010101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01000100010101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01000100010101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01000100010101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01000100010101010000) && ({row_reg, col_reg}<20'b01000100011000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01000100011000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01000100011000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01000100011000111000) && ({row_reg, col_reg}<20'b01000100011000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01000100011000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01000100011000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01000100011000111100) && ({row_reg, col_reg}<20'b01000100011000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01000100011000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01000100011000111111) && ({row_reg, col_reg}<20'b01000100011001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01000100011001100110) && ({row_reg, col_reg}<20'b01000100011001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01000100011001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01000100011001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01000100011001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01000100011001101011) && ({row_reg, col_reg}<20'b01000100100100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01000100100100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01000100100100011111) && ({row_reg, col_reg}<20'b01000100100101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01000100100101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01000100100101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01000100100101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01000100100101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01000100100101010000) && ({row_reg, col_reg}<20'b01000100101000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01000100101000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01000100101000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01000100101000111000) && ({row_reg, col_reg}<20'b01000100101000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01000100101000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01000100101000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01000100101000111100) && ({row_reg, col_reg}<20'b01000100101000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01000100101000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01000100101000111111) && ({row_reg, col_reg}<20'b01000100101001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01000100101001100110) && ({row_reg, col_reg}<20'b01000100101001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01000100101001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01000100101001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01000100101001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01000100101001101011) && ({row_reg, col_reg}<20'b01000100110100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01000100110100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01000100110100011111) && ({row_reg, col_reg}<20'b01000100110101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01000100110101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01000100110101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01000100110101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01000100110101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01000100110101010000) && ({row_reg, col_reg}<20'b01000100111000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01000100111000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01000100111000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01000100111000111000) && ({row_reg, col_reg}<20'b01000100111000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01000100111000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01000100111000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01000100111000111100) && ({row_reg, col_reg}<20'b01000100111000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01000100111000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01000100111000111111) && ({row_reg, col_reg}<20'b01000100111001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01000100111001100110) && ({row_reg, col_reg}<20'b01000100111001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01000100111001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01000100111001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01000100111001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01000100111001101011) && ({row_reg, col_reg}<20'b01000101000100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01000101000100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01000101000100011111) && ({row_reg, col_reg}<20'b01000101000101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01000101000101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01000101000101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01000101000101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01000101000101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01000101000101010000) && ({row_reg, col_reg}<20'b01000101001000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01000101001000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01000101001000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01000101001000111000) && ({row_reg, col_reg}<20'b01000101001000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01000101001000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01000101001000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01000101001000111100) && ({row_reg, col_reg}<20'b01000101001000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01000101001000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01000101001000111111) && ({row_reg, col_reg}<20'b01000101001001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01000101001001100110) && ({row_reg, col_reg}<20'b01000101001001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01000101001001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01000101001001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01000101001001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01000101001001101011) && ({row_reg, col_reg}<20'b01000101010100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01000101010100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01000101010100011111) && ({row_reg, col_reg}<20'b01000101010101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01000101010101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01000101010101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01000101010101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01000101010101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01000101010101010000) && ({row_reg, col_reg}<20'b01000101011000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01000101011000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01000101011000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01000101011000111000) && ({row_reg, col_reg}<20'b01000101011000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01000101011000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01000101011000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01000101011000111100) && ({row_reg, col_reg}<20'b01000101011000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01000101011000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01000101011000111111) && ({row_reg, col_reg}<20'b01000101011001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01000101011001100110) && ({row_reg, col_reg}<20'b01000101011001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01000101011001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01000101011001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01000101011001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01000101011001101011) && ({row_reg, col_reg}<20'b01000101100100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01000101100100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01000101100100011111) && ({row_reg, col_reg}<20'b01000101100101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01000101100101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01000101100101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01000101100101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01000101100101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01000101100101010000) && ({row_reg, col_reg}<20'b01000101101000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01000101101000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01000101101000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01000101101000111000) && ({row_reg, col_reg}<20'b01000101101000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01000101101000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01000101101000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01000101101000111100) && ({row_reg, col_reg}<20'b01000101101000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01000101101000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01000101101000111111) && ({row_reg, col_reg}<20'b01000101101001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01000101101001100110) && ({row_reg, col_reg}<20'b01000101101001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01000101101001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01000101101001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01000101101001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01000101101001101011) && ({row_reg, col_reg}<20'b01000101110100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01000101110100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01000101110100011111) && ({row_reg, col_reg}<20'b01000101110101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01000101110101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01000101110101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01000101110101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01000101110101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01000101110101010000) && ({row_reg, col_reg}<20'b01000101111000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01000101111000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01000101111000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01000101111000111000) && ({row_reg, col_reg}<20'b01000101111000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01000101111000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01000101111000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01000101111000111100) && ({row_reg, col_reg}<20'b01000101111000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01000101111000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01000101111000111111) && ({row_reg, col_reg}<20'b01000101111001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01000101111001100110) && ({row_reg, col_reg}<20'b01000101111001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01000101111001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01000101111001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01000101111001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01000101111001101011) && ({row_reg, col_reg}<20'b01000110000100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01000110000100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01000110000100011111) && ({row_reg, col_reg}<20'b01000110000101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01000110000101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01000110000101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01000110000101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01000110000101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01000110000101010000) && ({row_reg, col_reg}<20'b01000110001000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01000110001000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01000110001000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01000110001000111000) && ({row_reg, col_reg}<20'b01000110001000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01000110001000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01000110001000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01000110001000111100) && ({row_reg, col_reg}<20'b01000110001000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01000110001000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01000110001000111111) && ({row_reg, col_reg}<20'b01000110001001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01000110001001100110) && ({row_reg, col_reg}<20'b01000110001001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01000110001001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01000110001001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01000110001001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01000110001001101011) && ({row_reg, col_reg}<20'b01000110010100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01000110010100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01000110010100011111) && ({row_reg, col_reg}<20'b01000110010101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01000110010101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01000110010101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01000110010101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01000110010101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01000110010101010000) && ({row_reg, col_reg}<20'b01000110011000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01000110011000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01000110011000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01000110011000111000) && ({row_reg, col_reg}<20'b01000110011000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01000110011000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01000110011000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01000110011000111100) && ({row_reg, col_reg}<20'b01000110011000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01000110011000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01000110011000111111) && ({row_reg, col_reg}<20'b01000110011001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01000110011001100110) && ({row_reg, col_reg}<20'b01000110011001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01000110011001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01000110011001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01000110011001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01000110011001101011) && ({row_reg, col_reg}<20'b01000110100100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01000110100100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01000110100100011111) && ({row_reg, col_reg}<20'b01000110100101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01000110100101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01000110100101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01000110100101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01000110100101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01000110100101010000) && ({row_reg, col_reg}<20'b01000110101000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01000110101000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01000110101000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01000110101000111000) && ({row_reg, col_reg}<20'b01000110101000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01000110101000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01000110101000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01000110101000111100) && ({row_reg, col_reg}<20'b01000110101000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01000110101000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01000110101000111111) && ({row_reg, col_reg}<20'b01000110101001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01000110101001100110) && ({row_reg, col_reg}<20'b01000110101001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01000110101001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01000110101001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01000110101001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01000110101001101011) && ({row_reg, col_reg}<20'b01000110110100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01000110110100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01000110110100011111) && ({row_reg, col_reg}<20'b01000110110101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01000110110101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01000110110101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01000110110101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01000110110101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01000110110101010000) && ({row_reg, col_reg}<20'b01000110111000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01000110111000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01000110111000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01000110111000111000) && ({row_reg, col_reg}<20'b01000110111000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01000110111000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01000110111000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01000110111000111100) && ({row_reg, col_reg}<20'b01000110111000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01000110111000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01000110111000111111) && ({row_reg, col_reg}<20'b01000110111001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01000110111001100110) && ({row_reg, col_reg}<20'b01000110111001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01000110111001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01000110111001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01000110111001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01000110111001101011) && ({row_reg, col_reg}<20'b01000111000100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01000111000100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01000111000100011111) && ({row_reg, col_reg}<20'b01000111000101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01000111000101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01000111000101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01000111000101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01000111000101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01000111000101010000) && ({row_reg, col_reg}<20'b01000111001000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01000111001000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01000111001000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01000111001000111000) && ({row_reg, col_reg}<20'b01000111001000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01000111001000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01000111001000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01000111001000111100) && ({row_reg, col_reg}<20'b01000111001000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01000111001000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01000111001000111111) && ({row_reg, col_reg}<20'b01000111001001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01000111001001100110) && ({row_reg, col_reg}<20'b01000111001001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01000111001001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01000111001001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01000111001001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01000111001001101011) && ({row_reg, col_reg}<20'b01000111010100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01000111010100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01000111010100011111) && ({row_reg, col_reg}<20'b01000111010101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01000111010101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01000111010101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01000111010101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01000111010101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01000111010101010000) && ({row_reg, col_reg}<20'b01000111011000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01000111011000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01000111011000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01000111011000111000) && ({row_reg, col_reg}<20'b01000111011000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01000111011000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01000111011000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01000111011000111100) && ({row_reg, col_reg}<20'b01000111011000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01000111011000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01000111011000111111) && ({row_reg, col_reg}<20'b01000111011001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01000111011001100110) && ({row_reg, col_reg}<20'b01000111011001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01000111011001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01000111011001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01000111011001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01000111011001101011) && ({row_reg, col_reg}<20'b01000111100100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01000111100100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01000111100100011111) && ({row_reg, col_reg}<20'b01000111100101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01000111100101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01000111100101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01000111100101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01000111100101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01000111100101010000) && ({row_reg, col_reg}<20'b01000111101000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01000111101000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01000111101000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01000111101000111000) && ({row_reg, col_reg}<20'b01000111101000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01000111101000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01000111101000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01000111101000111100) && ({row_reg, col_reg}<20'b01000111101000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01000111101000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01000111101000111111) && ({row_reg, col_reg}<20'b01000111101001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01000111101001100110) && ({row_reg, col_reg}<20'b01000111101001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01000111101001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01000111101001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01000111101001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01000111101001101011) && ({row_reg, col_reg}<20'b01000111110100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01000111110100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01000111110100011111) && ({row_reg, col_reg}<20'b01000111110101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01000111110101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01000111110101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01000111110101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01000111110101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01000111110101010000) && ({row_reg, col_reg}<20'b01000111111000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01000111111000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01000111111000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01000111111000111000) && ({row_reg, col_reg}<20'b01000111111000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01000111111000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01000111111000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01000111111000111100) && ({row_reg, col_reg}<20'b01000111111000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01000111111000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01000111111000111111) && ({row_reg, col_reg}<20'b01000111111001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01000111111001100110) && ({row_reg, col_reg}<20'b01000111111001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01000111111001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01000111111001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01000111111001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01000111111001101011) && ({row_reg, col_reg}<20'b01001000000000001101)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=20'b01001000000000001101) && ({row_reg, col_reg}<20'b01001000000000001111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=20'b01001000000000001111) && ({row_reg, col_reg}<20'b01001000000000010110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01001000000000010110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=20'b01001000000000010111) && ({row_reg, col_reg}<20'b01001000000100011100)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01001000000100011100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==20'b01001000000100011101)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01001000000100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01001000000100011111) && ({row_reg, col_reg}<20'b01001000000101001001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01001000000101001001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01001000000101001010) && ({row_reg, col_reg}<20'b01001000000101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01001000000101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01001000000101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01001000000101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01001000000101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01001000000101010000) && ({row_reg, col_reg}<20'b01001000001000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01001000001000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01001000001000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01001000001000111000) && ({row_reg, col_reg}<20'b01001000001000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01001000001000111010) && ({row_reg, col_reg}<20'b01001000001000111111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01001000001000111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01001000001001000000) && ({row_reg, col_reg}<20'b01001000001001100000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01001000001001100000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01001000001001100001) && ({row_reg, col_reg}<20'b01001000001001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01001000001001100110) && ({row_reg, col_reg}<20'b01001000001001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01001000001001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01001000001001101001) && ({row_reg, col_reg}<20'b01001000001101110111)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01001000001101110111)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01001000001101111000) && ({row_reg, col_reg}<20'b01001000010000001010)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=20'b01001000010000001010) && ({row_reg, col_reg}<20'b01001000010000001100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=20'b01001000010000001100) && ({row_reg, col_reg}<20'b01001000010000010000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01001000010000010000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=20'b01001000010000010001) && ({row_reg, col_reg}<20'b01001000010000011010)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=20'b01001000010000011010) && ({row_reg, col_reg}<20'b01001000010100011110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01001000010100011110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==20'b01001000010100011111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01001000010100100000) && ({row_reg, col_reg}<20'b01001000010101001001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01001000010101001001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01001000010101001010) && ({row_reg, col_reg}<20'b01001000010101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01001000010101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01001000010101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01001000010101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01001000010101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==20'b01001000010101010000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=20'b01001000010101010001) && ({row_reg, col_reg}<20'b01001000011000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01001000011000110110)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==20'b01001000011000110111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=20'b01001000011000111000) && ({row_reg, col_reg}<20'b01001000011000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01001000011000111010) && ({row_reg, col_reg}<20'b01001000011001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01001000011001100110) && ({row_reg, col_reg}<20'b01001000011001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01001000011001101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01001000011001101001) && ({row_reg, col_reg}<20'b01001000011101101101)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=20'b01001000011101101101) && ({row_reg, col_reg}<20'b01001000011101110010)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01001000011101110010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=20'b01001000011101110011) && ({row_reg, col_reg}<20'b01001000011101111100)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=20'b01001000011101111100) && ({row_reg, col_reg}<20'b01001000011101111110)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01001000011101111110) && ({row_reg, col_reg}<20'b01001000100000001000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01001000100000001000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=20'b01001000100000001001) && ({row_reg, col_reg}<20'b01001000100000010110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=20'b01001000100000010110) && ({row_reg, col_reg}<20'b01001000100000011000)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=20'b01001000100000011000) && ({row_reg, col_reg}<20'b01001000100000011010)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=20'b01001000100000011010) && ({row_reg, col_reg}<20'b01001000100000011100)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01001000100000011100) && ({row_reg, col_reg}<20'b01001000100100011110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==20'b01001000100100011110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=20'b01001000100100011111) && ({row_reg, col_reg}<20'b01001000100101001001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01001000100101001001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01001000100101001010) && ({row_reg, col_reg}<20'b01001000100101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01001000100101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01001000100101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01001000100101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01001000100101001111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=20'b01001000100101010000) && ({row_reg, col_reg}<20'b01001000101000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01001000101000110111) && ({row_reg, col_reg}<20'b01001000101000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01001000101000111010) && ({row_reg, col_reg}<20'b01001000101000111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01001000101000111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01001000101000111101) && ({row_reg, col_reg}<20'b01001000101001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01001000101001100110) && ({row_reg, col_reg}<20'b01001000101001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01001000101001101000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=20'b01001000101001101001) && ({row_reg, col_reg}<20'b01001000101101101011)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01001000101101101011) && ({row_reg, col_reg}<20'b01001000101101101101)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01001000101101101101) && ({row_reg, col_reg}<20'b01001000101101101111)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=20'b01001000101101101111) && ({row_reg, col_reg}<20'b01001000101101110001)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=20'b01001000101101110001) && ({row_reg, col_reg}<20'b01001000101101110101)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=20'b01001000101101110101) && ({row_reg, col_reg}<20'b01001000101101110111)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01001000101101110111) && ({row_reg, col_reg}<20'b01001000110000001100)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=20'b01001000110000001100) && ({row_reg, col_reg}<20'b01001000110000001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=20'b01001000110000001110) && ({row_reg, col_reg}<20'b01001000110000010010)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01001000110000010010)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01001000110000010011)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==20'b01001000110000010100)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01001000110000010101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01001000110000010110) && ({row_reg, col_reg}<20'b01001000110000011001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=20'b01001000110000011001) && ({row_reg, col_reg}<20'b01001000110100011111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01001000110100011111) && ({row_reg, col_reg}<20'b01001000110101001001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01001000110101001001) && ({row_reg, col_reg}<20'b01001000110101001011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01001000110101001011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01001000110101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01001000110101001101) && ({row_reg, col_reg}<20'b01001000110101001111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01001000110101001111) && ({row_reg, col_reg}<20'b01001000111000111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01001000111000111001) && ({row_reg, col_reg}<20'b01001000111000111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01001000111000111100) && ({row_reg, col_reg}<20'b01001000111000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01001000111000111110) && ({row_reg, col_reg}<20'b01001000111001100111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01001000111001100111) && ({row_reg, col_reg}<20'b01001000111101101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01001000111101101110) && ({row_reg, col_reg}<20'b01001000111101110001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==20'b01001000111101110001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==20'b01001000111101110010)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01001000111101110011)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==20'b01001000111101110100)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01001000111101110101)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=20'b01001000111101110110) && ({row_reg, col_reg}<20'b01001000111101111000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=20'b01001000111101111000) && ({row_reg, col_reg}<20'b01001000111101111010)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01001000111101111010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=20'b01001000111101111011) && ({row_reg, col_reg}<20'b01001000111101111110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=20'b01001000111101111110) && ({row_reg, col_reg}<20'b01001000111110000000)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01001000111110000000) && ({row_reg, col_reg}<20'b01001001000000010000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01001001000000010000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==20'b01001001000000010001)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01001001000000010010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01001001000000010011) && ({row_reg, col_reg}<20'b01001001000000010101)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=20'b01001001000000010101) && ({row_reg, col_reg}<20'b01001001000000011000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01001001000000011000) && ({row_reg, col_reg}<20'b01001001000000011010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01001001000000011010) && ({row_reg, col_reg}<20'b01001001000000100000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01001001000000100000) && ({row_reg, col_reg}<20'b01001001000100011100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01001001000100011100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01001001000100011101) && ({row_reg, col_reg}<20'b01001001000100011111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01001001000100011111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01001001000100100000) && ({row_reg, col_reg}<20'b01001001000101001001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01001001000101001001) && ({row_reg, col_reg}<20'b01001001000101001011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01001001000101001011) && ({row_reg, col_reg}<20'b01001001000101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01001001000101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01001001000101010010) && ({row_reg, col_reg}<20'b01001001001000110011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01001001001000110011) && ({row_reg, col_reg}<20'b01001001001000110101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01001001001000110101) && ({row_reg, col_reg}<20'b01001001001000110111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01001001001000110111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01001001001000111000) && ({row_reg, col_reg}<20'b01001001001000111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01001001001000111101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01001001001000111110) && ({row_reg, col_reg}<20'b01001001001001101110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01001001001001101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01001001001001101111) && ({row_reg, col_reg}<20'b01001001001101101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01001001001101101000) && ({row_reg, col_reg}<20'b01001001001101101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01001001001101101100) && ({row_reg, col_reg}<20'b01001001001101110000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01001001001101110000) && ({row_reg, col_reg}<20'b01001001001101110011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01001001001101110011)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==20'b01001001001101110100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==20'b01001001001101110101)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01001001001101110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=20'b01001001001101110111) && ({row_reg, col_reg}<20'b01001001001101111101)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=20'b01001001001101111101) && ({row_reg, col_reg}<20'b01001001001101111111)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01001001001101111111) && ({row_reg, col_reg}<20'b01001001010000001001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01001001010000001001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=20'b01001001010000001010) && ({row_reg, col_reg}<20'b01001001010000001110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01001001010000001110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01001001010000001111)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==20'b01001001010000010000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==20'b01001001010000010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01001001010000010010) && ({row_reg, col_reg}<20'b01001001010000011010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01001001010000011010) && ({row_reg, col_reg}<20'b01001001010000011100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01001001010000011100) && ({row_reg, col_reg}<20'b01001001010000100000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01001001010000100000) && ({row_reg, col_reg}<20'b01001001010100011001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01001001010100011001) && ({row_reg, col_reg}<20'b01001001010100011011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01001001010100011011) && ({row_reg, col_reg}<20'b01001001010100011101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01001001010100011101) && ({row_reg, col_reg}<20'b01001001010101001001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01001001010101001001) && ({row_reg, col_reg}<20'b01001001010101001011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01001001010101001011) && ({row_reg, col_reg}<20'b01001001010101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01001001010101001101) && ({row_reg, col_reg}<20'b01001001010101001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01001001010101001111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01001001010101010000) && ({row_reg, col_reg}<20'b01001001010101010010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01001001010101010010) && ({row_reg, col_reg}<20'b01001001010101010100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01001001010101010100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01001001010101010101) && ({row_reg, col_reg}<20'b01001001010101010111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01001001010101010111) && ({row_reg, col_reg}<20'b01001001011000110001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01001001011000110001) && ({row_reg, col_reg}<20'b01001001011000110100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01001001011000110100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01001001011000110101) && ({row_reg, col_reg}<20'b01001001011000110111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01001001011000110111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01001001011000111000) && ({row_reg, col_reg}<20'b01001001011000111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01001001011000111101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01001001011000111110) && ({row_reg, col_reg}<20'b01001001011001100010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01001001011001100010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01001001011001100011) && ({row_reg, col_reg}<20'b01001001011001101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01001001011001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01001001011001101001) && ({row_reg, col_reg}<20'b01001001011001101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01001001011001101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01001001011001101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01001001011001101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01001001011001101111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01001001011001110000) && ({row_reg, col_reg}<20'b01001001011101101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01001001011101101000) && ({row_reg, col_reg}<20'b01001001011101101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01001001011101101101) && ({row_reg, col_reg}<20'b01001001011101110000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01001001011101110000) && ({row_reg, col_reg}<20'b01001001011101110100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01001001011101110100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01001001011101110101)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==20'b01001001011101110110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01001001011101110111)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=20'b01001001011101111000) && ({row_reg, col_reg}<20'b01001001011101111010)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=20'b01001001011101111010) && ({row_reg, col_reg}<20'b01001001011101111100)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01001001011101111100) && ({row_reg, col_reg}<20'b01001001100000001101)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01001001100000001101)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01001001100000001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01001001100000001111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==20'b01001001100000010000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01001001100000010001) && ({row_reg, col_reg}<20'b01001001100000010100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01001001100000010100) && ({row_reg, col_reg}<20'b01001001100000011000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01001001100000011000) && ({row_reg, col_reg}<20'b01001001100000011111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01001001100000011111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01001001100000100000) && ({row_reg, col_reg}<20'b01001001100100011001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01001001100100011001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01001001100100011010) && ({row_reg, col_reg}<20'b01001001100101001010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01001001100101001010) && ({row_reg, col_reg}<20'b01001001100101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01001001100101001100) && ({row_reg, col_reg}<20'b01001001100101001110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01001001100101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01001001100101001111) && ({row_reg, col_reg}<20'b01001001100101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01001001100101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01001001100101010010) && ({row_reg, col_reg}<20'b01001001100101010100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01001001100101010100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01001001100101010101) && ({row_reg, col_reg}<20'b01001001100101010111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01001001100101010111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01001001100101011000) && ({row_reg, col_reg}<20'b01001001101000110000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01001001101000110000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01001001101000110001) && ({row_reg, col_reg}<20'b01001001101000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01001001101000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01001001101000111011) && ({row_reg, col_reg}<20'b01001001101000111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01001001101000111101) && ({row_reg, col_reg}<20'b01001001101000111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01001001101000111111) && ({row_reg, col_reg}<20'b01001001101001100001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01001001101001100001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01001001101001100010) && ({row_reg, col_reg}<20'b01001001101001100101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01001001101001100101) && ({row_reg, col_reg}<20'b01001001101001100111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01001001101001100111) && ({row_reg, col_reg}<20'b01001001101001101010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01001001101001101010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01001001101001101011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01001001101001101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01001001101001101101) && ({row_reg, col_reg}<20'b01001001101001101111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01001001101001101111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01001001101001110000) && ({row_reg, col_reg}<20'b01001001101101101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01001001101101101000) && ({row_reg, col_reg}<20'b01001001101101101011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01001001101101101011) && ({row_reg, col_reg}<20'b01001001101101110001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01001001101101110001) && ({row_reg, col_reg}<20'b01001001101101110100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01001001101101110100) && ({row_reg, col_reg}<20'b01001001101101110110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01001001101101110110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01001001101101110111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==20'b01001001101101111000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01001001101101111001)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01001001101101111010)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01001001101101111011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=20'b01001001101101111100) && ({row_reg, col_reg}<20'b01001001101101111111)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01001001101101111111)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01001001101110000000) && ({row_reg, col_reg}<20'b01001001110000001011)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01001001110000001011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01001001110000001100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==20'b01001001110000001101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01001001110000001110) && ({row_reg, col_reg}<20'b01001001110000010000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01001001110000010000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01001001110000010001) && ({row_reg, col_reg}<20'b01001001110000010011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01001001110000010011) && ({row_reg, col_reg}<20'b01001001110000010110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01001001110000010110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01001001110000010111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01001001110000011000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01001001110000011001) && ({row_reg, col_reg}<20'b01001001110000011101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01001001110000011101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01001001110000011110) && ({row_reg, col_reg}<20'b01001001110100011001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01001001110100011001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01001001110100011010) && ({row_reg, col_reg}<20'b01001001110100011101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01001001110100011101) && ({row_reg, col_reg}<20'b01001001110100011111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01001001110100011111) && ({row_reg, col_reg}<20'b01001001110101001010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01001001110101001010) && ({row_reg, col_reg}<20'b01001001110101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01001001110101001100) && ({row_reg, col_reg}<20'b01001001110101001110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01001001110101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01001001110101001111) && ({row_reg, col_reg}<20'b01001001110101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01001001110101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01001001110101010010) && ({row_reg, col_reg}<20'b01001001110101010100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01001001110101010100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01001001110101010101) && ({row_reg, col_reg}<20'b01001001110101010111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01001001110101010111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01001001110101011000) && ({row_reg, col_reg}<20'b01001001111000110000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01001001111000110000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01001001111000110001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01001001111000110010) && ({row_reg, col_reg}<20'b01001001111000110100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01001001111000110100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01001001111000110101) && ({row_reg, col_reg}<20'b01001001111000110111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01001001111000110111) && ({row_reg, col_reg}<20'b01001001111000111001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01001001111000111001) && ({row_reg, col_reg}<20'b01001001111000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01001001111000111011) && ({row_reg, col_reg}<20'b01001001111000111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01001001111000111101) && ({row_reg, col_reg}<20'b01001001111000111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01001001111000111111) && ({row_reg, col_reg}<20'b01001001111001100001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01001001111001100001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01001001111001100010) && ({row_reg, col_reg}<20'b01001001111001100101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01001001111001100101) && ({row_reg, col_reg}<20'b01001001111001100111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01001001111001100111) && ({row_reg, col_reg}<20'b01001001111001101010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01001001111001101010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01001001111001101011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01001001111001101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01001001111001101101) && ({row_reg, col_reg}<20'b01001001111001101111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01001001111001101111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01001001111001110000) && ({row_reg, col_reg}<20'b01001001111101110000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01001001111101110000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01001001111101110001) && ({row_reg, col_reg}<20'b01001001111101110011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01001001111101110011) && ({row_reg, col_reg}<20'b01001001111101111000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01001001111101111000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==20'b01001001111101111001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==20'b01001001111101111010)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==20'b01001001111101111011)) color_data = 12'b110111011101;

		if(({row_reg, col_reg}>=20'b01001001111101111100) && ({row_reg, col_reg}<20'b01001010000000000000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01001010000000000000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==20'b01001010000000000001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01001010000000000010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=20'b01001010000000000011) && ({row_reg, col_reg}<20'b01001010000000001010)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01001010000000001010)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01001010000000001011)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01001010000000001100)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==20'b01001010000000001101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01001010000000001110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01001010000000001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01001010000000010000) && ({row_reg, col_reg}<20'b01001010001101111001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01001010001101111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01001010001101111010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==20'b01001010001101111011)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01001010001101111100)) color_data = 12'b110111011101;

		if(({row_reg, col_reg}>=20'b01001010001101111101) && ({row_reg, col_reg}<20'b01001010010000000111)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01001010010000000111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==20'b01001010010000001000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01001010010000001001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==20'b01001010010000001010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==20'b01001010010000001011)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==20'b01001010010000001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01001010010000001101) && ({row_reg, col_reg}<20'b01001010011101111000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01001010011101111000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01001010011101111001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01001010011101111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01001010011101111011)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==20'b01001010011101111100)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01001010011101111101)) color_data = 12'b110111011101;

		if(({row_reg, col_reg}>=20'b01001010011101111110) && ({row_reg, col_reg}<20'b01001010100000000001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01001010100000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=20'b01001010100000000010) && ({row_reg, col_reg}<20'b01001010100000001000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01001010100000001000)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01001010100000001001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==20'b01001010100000001010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01001010100000001011) && ({row_reg, col_reg}<20'b01001010100000001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01001010100000001101) && ({row_reg, col_reg}<20'b01001010100000010000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01001010100000010000) && ({row_reg, col_reg}<20'b01001010101101111000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01001010101101111000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01001010101101111001) && ({row_reg, col_reg}<20'b01001010101101111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01001010101101111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01001010101101111101)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01001010101101111110) && ({row_reg, col_reg}<20'b01001010101110000010)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01001010101110000010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01001010101110000011) && ({row_reg, col_reg}<20'b01001010110000000001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01001010110000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=20'b01001010110000000010) && ({row_reg, col_reg}<20'b01001010110000000101)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=20'b01001010110000000101) && ({row_reg, col_reg}<20'b01001010110000000111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==20'b01001010110000000111)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01001010110000001000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01001010110000001001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==20'b01001010110000001010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01001010110000001011) && ({row_reg, col_reg}<20'b01001010110000001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01001010110000001110) && ({row_reg, col_reg}<20'b01001010111101111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01001010111101111010) && ({row_reg, col_reg}<20'b01001010111101111101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01001010111101111101)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==20'b01001010111101111110)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=20'b01001010111101111111) && ({row_reg, col_reg}<20'b01001010111110000011)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}==20'b01001010111110000011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=20'b01001011000000000000) && ({row_reg, col_reg}<20'b01001011000000000101)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01001011000000000101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==20'b01001011000000000110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01001011000000000111)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==20'b01001011000000001000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==20'b01001011000000001001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01001011000000001010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01001011000000001011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01001011000000001100) && ({row_reg, col_reg}<20'b01001011000000001111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01001011000000001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01001011000000010000) && ({row_reg, col_reg}<20'b01001011001101111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01001011001101111100) && ({row_reg, col_reg}<20'b01001011001101111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01001011001101111110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==20'b01001011001101111111)) color_data = 12'b110111011101;

		if(({row_reg, col_reg}>=20'b01001011001110000000) && ({row_reg, col_reg}<20'b01001011010000000011)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01001011010000000011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=20'b01001011010000000100) && ({row_reg, col_reg}<20'b01001011010000000110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01001011010000000110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01001011010000000111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==20'b01001011010000001000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01001011010000001001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01001011010000001010) && ({row_reg, col_reg}<20'b01001011010000001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01001011010000001100) && ({row_reg, col_reg}<20'b01001011010000001110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01001011010000001110) && ({row_reg, col_reg}<20'b01001011010000010000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01001011010000010000) && ({row_reg, col_reg}<20'b01001011011101111001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01001011011101111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01001011011101111010) && ({row_reg, col_reg}<20'b01001011011101111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01001011011101111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01001011011101111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01001011011101111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01001011011101111111)) color_data = 12'b101110111011;

		if(({row_reg, col_reg}>=20'b01001011011110000000) && ({row_reg, col_reg}<20'b01001011100000000000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01001011100000000000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==20'b01001011100000000001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01001011100000000010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=20'b01001011100000000011) && ({row_reg, col_reg}<20'b01001011100000000110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01001011100000000110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01001011100000000111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=20'b01001011100000001000) && ({row_reg, col_reg}<20'b01001011100000001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01001011100000001101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01001011100000001110) && ({row_reg, col_reg}<20'b01001011101101111001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01001011101101111001) && ({row_reg, col_reg}<20'b01001011101101111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01001011101101111011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01001011101101111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01001011101101111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01001011101101111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01001011101101111111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==20'b01001011101110000000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==20'b01001011101110000001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01001011101110000010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01001011101110000011) && ({row_reg, col_reg}<20'b01001011110000000101)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01001011110000000101)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01001011110000000110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=20'b01001011110000000111) && ({row_reg, col_reg}<20'b01001011110000001011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01001011110000001011) && ({row_reg, col_reg}<20'b01001011110000001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01001011110000001101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01001011110000001110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01001011110000001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01001011110000010000) && ({row_reg, col_reg}<20'b01001011111101111011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01001011111101111011) && ({row_reg, col_reg}<20'b01001011111101111101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01001011111101111101) && ({row_reg, col_reg}<20'b01001011111101111111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01001011111101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01001011111110000000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==20'b01001011111110000001)) color_data = 12'b110111011101;

		if(({row_reg, col_reg}>=20'b01001011111110000010) && ({row_reg, col_reg}<20'b01001100000000000000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01001100000000000000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=20'b01001100000000000001) && ({row_reg, col_reg}<20'b01001100000000000011)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01001100000000000011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==20'b01001100000000000100)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01001100000000000101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01001100000000000110) && ({row_reg, col_reg}<20'b01001100000000001000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01001100000000001000) && ({row_reg, col_reg}<20'b01001100001110000000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01001100001110000000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01001100001110000001)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01001100001110000010)) color_data = 12'b110111011101;

		if(({row_reg, col_reg}>=20'b01001100001110000011) && ({row_reg, col_reg}<20'b01001100010000000100)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01001100010000000100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==20'b01001100010000000101)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==20'b01001100010000000110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01001100010000000111) && ({row_reg, col_reg}<20'b01001100011110000000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01001100011110000000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01001100011110000001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==20'b01001100011110000010)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=20'b01001100011110000011) && ({row_reg, col_reg}<20'b01001100100000000001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01001100100000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=20'b01001100100000000010) && ({row_reg, col_reg}<20'b01001100100000000100)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01001100100000000100)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01001100100000000101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01001100100000000110) && ({row_reg, col_reg}<20'b01001100101110000000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01001100101110000000) && ({row_reg, col_reg}<20'b01001100101110000010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01001100101110000010)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=20'b01001100101110000011) && ({row_reg, col_reg}<20'b01001100110000000001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01001100110000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==20'b01001100110000000010)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01001100110000000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01001100110000000100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==20'b01001100110000000101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01001100110000000110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01001100110000000111) && ({row_reg, col_reg}<20'b01001100111110000000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01001100111110000000) && ({row_reg, col_reg}<20'b01001100111110000010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01001100111110000010)) color_data = 12'b101110111011;

		if(({row_reg, col_reg}>=20'b01001100111110000011) && ({row_reg, col_reg}<20'b01001101000000000011)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01001101000000000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01001101000000000100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==20'b01001101000000000101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01001101000000000110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01001101000000000111) && ({row_reg, col_reg}<20'b01001101001110000010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01001101001110000010)) color_data = 12'b101110111011;

		if(({row_reg, col_reg}>=20'b01001101001110000011) && ({row_reg, col_reg}<20'b01001101010000000011)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01001101010000000011)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==20'b01001101010000000100)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==20'b01001101010000000101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01001101010000000110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01001101010000000111) && ({row_reg, col_reg}<20'b01001101011110000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01001101011110000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01001101011110000010)) color_data = 12'b101010101010;

		if(({row_reg, col_reg}==20'b01001101011110000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=20'b01001101100000000000) && ({row_reg, col_reg}<20'b01001101100000000011)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01001101100000000011)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01001101100000000100)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=20'b01001101100000000101) && ({row_reg, col_reg}<20'b01001101100000000111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01001101100000000111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01001101100000001000) && ({row_reg, col_reg}<20'b01001101101110000000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01001101101110000000) && ({row_reg, col_reg}<20'b01001101101110000010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01001101101110000010)) color_data = 12'b100110011001;

		if(({row_reg, col_reg}==20'b01001101101110000011)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01001101110000000000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=20'b01001101110000000001) && ({row_reg, col_reg}<20'b01001101110000000011)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01001101110000000011)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01001101110000000100) && ({row_reg, col_reg}<20'b01001101110000000110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01001101110000000110) && ({row_reg, col_reg}<20'b01001101111110000010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01001101111110000010)) color_data = 12'b100110011001;

		if(({row_reg, col_reg}==20'b01001101111110000011)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01001110000000000000) && ({row_reg, col_reg}<20'b01001110000000000011)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01001110000000000011)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01001110000000000100) && ({row_reg, col_reg}<20'b01001110000000000110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01001110000000000110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01001110000000000111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01001110000000001000) && ({row_reg, col_reg}<20'b01001110001110000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01001110001110000001) && ({row_reg, col_reg}<20'b01001110001110000011)) color_data = 12'b100010001000;

		if(({row_reg, col_reg}==20'b01001110001110000011)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=20'b01001110010000000000) && ({row_reg, col_reg}<20'b01001110010000000010)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01001110010000000010)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01001110010000000011)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=20'b01001110010000000100) && ({row_reg, col_reg}<20'b01001110010000000110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01001110010000000110) && ({row_reg, col_reg}<20'b01001110011110000010)) color_data = 12'b011101110111;

		if(({row_reg, col_reg}>=20'b01001110011110000010) && ({row_reg, col_reg}<20'b01001110100000000000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01001110100000000000) && ({row_reg, col_reg}<20'b01001110100000000010)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01001110100000000010)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01001110100000000011)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=20'b01001110100000000100) && ({row_reg, col_reg}<20'b01001110101110000000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01001110101110000000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01001110101110000001)) color_data = 12'b011101110111;

		if(({row_reg, col_reg}>=20'b01001110101110000010) && ({row_reg, col_reg}<20'b01001110110000000000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01001110110000000000) && ({row_reg, col_reg}<20'b01001110110000000010)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01001110110000000010)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01001110110000000011)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=20'b01001110110000000100) && ({row_reg, col_reg}<20'b01001110110000000111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01001110110000000111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01001110110000001000) && ({row_reg, col_reg}<20'b01001110111110000000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01001110111110000000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01001110111110000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01001110111110000010)) color_data = 12'b100010001000;

		if(({row_reg, col_reg}==20'b01001110111110000011)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=20'b01001111000000000000) && ({row_reg, col_reg}<20'b01001111000000000010)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01001111000000000010)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01001111000000000011)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==20'b01001111000000000100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01001111000000000101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01001111000000000110) && ({row_reg, col_reg}<20'b01001111000000001000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01001111000000001000) && ({row_reg, col_reg}<20'b01001111001110000000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01001111001110000000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01001111001110000001)) color_data = 12'b011101110111;

		if(({row_reg, col_reg}>=20'b01001111001110000010) && ({row_reg, col_reg}<20'b01001111010000000000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=20'b01001111010000000000) && ({row_reg, col_reg}<20'b01001111010000000010)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01001111010000000010)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01001111010000000011)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==20'b01001111010000000100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01001111010000000101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01001111010000000110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01001111010000000111) && ({row_reg, col_reg}<20'b01001111011110000000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01001111011110000000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01001111011110000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01001111011110000010)) color_data = 12'b100110011001;

		if(({row_reg, col_reg}==20'b01001111011110000011)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01001111100000000000) && ({row_reg, col_reg}<20'b01001111100000000011)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01001111100000000011)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01001111100000000100)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==20'b01001111100000000101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01001111100000000110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01001111100000000111) && ({row_reg, col_reg}<20'b01001111101110000000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01001111101110000000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01001111101110000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01001111101110000010)) color_data = 12'b100110011001;

		if(({row_reg, col_reg}==20'b01001111101110000011)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01001111110000000000) && ({row_reg, col_reg}<20'b01001111110000000011)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01001111110000000011)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01001111110000000100)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==20'b01001111110000000101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01001111110000000110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01001111110000000111) && ({row_reg, col_reg}<20'b01001111111110000010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01001111111110000010)) color_data = 12'b101010101010;

		if(({row_reg, col_reg}==20'b01001111111110000011)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==20'b01010000000000000000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01010000000000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==20'b01010000000000000010)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01010000000000000011)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==20'b01010000000000000100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==20'b01010000000000000101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01010000000000000110) && ({row_reg, col_reg}<20'b01010000001101111001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01010000001101111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01010000001101111010) && ({row_reg, col_reg}<20'b01010000001101111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01010000001101111101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01010000001101111110) && ({row_reg, col_reg}<20'b01010000001110000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01010000001110000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01010000001110000010)) color_data = 12'b101010101010;

		if(({row_reg, col_reg}==20'b01010000001110000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01010000010000000000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01010000010000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==20'b01010000010000000010)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01010000010000000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01010000010000000100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==20'b01010000010000000101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01010000010000000110) && ({row_reg, col_reg}<20'b01010000010000001000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01010000010000001000) && ({row_reg, col_reg}<20'b01010000011101111011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01010000011101111011) && ({row_reg, col_reg}<20'b01010000011101111101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01010000011101111101) && ({row_reg, col_reg}<20'b01010000011110000010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01010000011110000010)) color_data = 12'b101110111011;

		if(({row_reg, col_reg}>=20'b01010000011110000011) && ({row_reg, col_reg}<20'b01010000100000000100)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01010000100000000100)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01010000100000000101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01010000100000000110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01010000100000000111) && ({row_reg, col_reg}<20'b01010000101101111000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01010000101101111000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01010000101101111001) && ({row_reg, col_reg}<20'b01010000101101111011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01010000101101111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01010000101101111100) && ({row_reg, col_reg}<20'b01010000101101111111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01010000101101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01010000101110000000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01010000101110000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01010000101110000010)) color_data = 12'b101110111011;

		if(({row_reg, col_reg}>=20'b01010000101110000011) && ({row_reg, col_reg}<20'b01010000110000000100)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01010000110000000100)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01010000110000000101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01010000110000000110) && ({row_reg, col_reg}<20'b01010000111101111000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01010000111101111000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01010000111101111001) && ({row_reg, col_reg}<20'b01010000111101111011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01010000111101111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01010000111101111100) && ({row_reg, col_reg}<20'b01010000111101111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01010000111101111110) && ({row_reg, col_reg}<20'b01010000111110000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01010000111110000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==20'b01010000111110000010)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}==20'b01010000111110000011)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01010001000000000000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=20'b01010001000000000001) && ({row_reg, col_reg}<20'b01010001000000000100)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01010001000000000100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==20'b01010001000000000101)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=20'b01010001000000000110) && ({row_reg, col_reg}<20'b01010001000000001000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01010001000000001000) && ({row_reg, col_reg}<20'b01010001001101111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01010001001101111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01010001001101111111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01010001001110000000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01010001001110000001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==20'b01010001001110000010)) color_data = 12'b110111011101;

		if(({row_reg, col_reg}>=20'b01010001001110000011) && ({row_reg, col_reg}<20'b01010001010000000010)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01010001010000000010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==20'b01010001010000000011)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01010001010000000100)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01010001010000000101)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01010001010000000110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01010001010000000111) && ({row_reg, col_reg}<20'b01010001011101111001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01010001011101111001) && ({row_reg, col_reg}<20'b01010001011101111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01010001011101111011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01010001011101111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01010001011101111101) && ({row_reg, col_reg}<20'b01010001011101111111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01010001011101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01010001011110000000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==20'b01010001011110000001)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=20'b01010001011110000010) && ({row_reg, col_reg}<20'b01010001100000000010)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01010001100000000010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=20'b01010001100000000011) && ({row_reg, col_reg}<20'b01010001100000000101)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01010001100000000101)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01010001100000000110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==20'b01010001100000000111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01010001100000001000) && ({row_reg, col_reg}<20'b01010001101101111001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01010001101101111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01010001101101111010) && ({row_reg, col_reg}<20'b01010001101101111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01010001101101111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01010001101101111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01010001101101111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01010001101101111111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==20'b01010001101110000000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01010001101110000001) && ({row_reg, col_reg}<20'b01010001101110000011)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}>=20'b01010001101110000011) && ({row_reg, col_reg}<20'b01010001110000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=20'b01010001110000000001) && ({row_reg, col_reg}<20'b01010001110000000100)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01010001110000000100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==20'b01010001110000000101)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01010001110000000110)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==20'b01010001110000000111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=20'b01010001110000001000) && ({row_reg, col_reg}<20'b01010001111101111001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01010001111101111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01010001111101111010) && ({row_reg, col_reg}<20'b01010001111101111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01010001111101111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01010001111101111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01010001111101111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01010001111101111111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==20'b01010001111110000000)) color_data = 12'b110111011101;

		if(({row_reg, col_reg}>=20'b01010001111110000001) && ({row_reg, col_reg}<20'b01010010000000000010)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01010010000000000010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=20'b01010010000000000011) && ({row_reg, col_reg}<20'b01010010000000000101)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01010010000000000101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==20'b01010010000000000110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01010010000000000111)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01010010000000001000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=20'b01010010000000001001) && ({row_reg, col_reg}<20'b01010010000000001011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01010010000000001011) && ({row_reg, col_reg}<20'b01010010000000001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01010010000000001101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01010010000000001110) && ({row_reg, col_reg}<20'b01010010000000010111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01010010000000010111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01010010000000011000) && ({row_reg, col_reg}<20'b01010010001101110000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01010010001101110000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01010010001101110001) && ({row_reg, col_reg}<20'b01010010001101110011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01010010001101110011) && ({row_reg, col_reg}<20'b01010010001101110101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01010010001101110101) && ({row_reg, col_reg}<20'b01010010001101111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01010010001101111010) && ({row_reg, col_reg}<20'b01010010001101111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01010010001101111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01010010001101111101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01010010001101111110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==20'b01010010001101111111)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=20'b01010010001110000000) && ({row_reg, col_reg}<20'b01010010010000000000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01010010010000000000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==20'b01010010010000000001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=20'b01010010010000000010) && ({row_reg, col_reg}<20'b01010010010000000100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==20'b01010010010000000100)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01010010010000000101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==20'b01010010010000000110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01010010010000000111)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01010010010000001000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01010010010000001001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01010010010000001010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01010010010000001011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01010010010000001100) && ({row_reg, col_reg}<20'b01010010010000001110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01010010010000001110) && ({row_reg, col_reg}<20'b01010010010000010110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01010010010000010110) && ({row_reg, col_reg}<20'b01010010011101110011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01010010011101110011) && ({row_reg, col_reg}<20'b01010010011101110110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01010010011101110110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01010010011101110111) && ({row_reg, col_reg}<20'b01010010011101111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01010010011101111010) && ({row_reg, col_reg}<20'b01010010011101111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01010010011101111101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01010010011101111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01010010011101111111)) color_data = 12'b110111011101;

		if(({row_reg, col_reg}>=20'b01010010011110000000) && ({row_reg, col_reg}<20'b01010010100000000000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01010010100000000000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=20'b01010010100000000001) && ({row_reg, col_reg}<20'b01010010100000000101)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=20'b01010010100000000101) && ({row_reg, col_reg}<20'b01010010100000000111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==20'b01010010100000000111)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01010010100000001000)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01010010100000001001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=20'b01010010100000001010) && ({row_reg, col_reg}<20'b01010010100000001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01010010100000001100) && ({row_reg, col_reg}<20'b01010010100000010100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01010010100000010100) && ({row_reg, col_reg}<20'b01010010100000010110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01010010100000010110) && ({row_reg, col_reg}<20'b01010010101101111001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01010010101101111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01010010101101111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01010010101101111011) && ({row_reg, col_reg}<20'b01010010101101111101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01010010101101111101)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==20'b01010010101101111110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01010010101101111111)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01010010101110000000) && ({row_reg, col_reg}<20'b01010010110000000111)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01010010110000000111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==20'b01010010110000001000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01010010110000001001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==20'b01010010110000001010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==20'b01010010110000001011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01010010110000001100) && ({row_reg, col_reg}<20'b01010010110000001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01010010110000001110) && ({row_reg, col_reg}<20'b01010010110000010110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01010010110000010110) && ({row_reg, col_reg}<20'b01010010110000011000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01010010110000011000) && ({row_reg, col_reg}<20'b01010010111101110110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01010010111101110110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01010010111101110111) && ({row_reg, col_reg}<20'b01010010111101111001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01010010111101111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01010010111101111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01010010111101111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01010010111101111100)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==20'b01010010111101111101)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=20'b01010010111101111110) && ({row_reg, col_reg}<20'b01010011000000000001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01010011000000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=20'b01010011000000000010) && ({row_reg, col_reg}<20'b01010011000000001010)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01010011000000001010)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01010011000000001011)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=20'b01010011000000001100) && ({row_reg, col_reg}<20'b01010011000000001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01010011000000001110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01010011000000001111) && ({row_reg, col_reg}<20'b01010011000000010011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01010011000000010011) && ({row_reg, col_reg}<20'b01010011000000010111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01010011000000010111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01010011000000011000) && ({row_reg, col_reg}<20'b01010011001101110101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01010011001101110101) && ({row_reg, col_reg}<20'b01010011001101110111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01010011001101110111) && ({row_reg, col_reg}<20'b01010011001101111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01010011001101111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01010011001101111011)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==20'b01010011001101111100)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01010011001101111101)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01010011001101111110)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01010011001101111111) && ({row_reg, col_reg}<20'b01010011010000000001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01010011010000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=20'b01010011010000000010) && ({row_reg, col_reg}<20'b01010011010000001010)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01010011010000001010)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01010011010000001011)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==20'b01010011010000001100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01010011010000001101) && ({row_reg, col_reg}<20'b01010011010000001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01010011010000001111) && ({row_reg, col_reg}<20'b01010011010000010011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01010011010000010011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01010011010000010100) && ({row_reg, col_reg}<20'b01010011011101110011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01010011011101110011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01010011011101110100) && ({row_reg, col_reg}<20'b01010011011101111000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01010011011101111000) && ({row_reg, col_reg}<20'b01010011011101111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01010011011101111010)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01010011011101111011)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==20'b01010011011101111100)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01010011011101111101)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01010011011101111110) && ({row_reg, col_reg}<20'b01010011100000001100)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01010011100000001100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==20'b01010011100000001101)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01010011100000001110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01010011100000001111) && ({row_reg, col_reg}<20'b01010011100000010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01010011100000010001) && ({row_reg, col_reg}<20'b01010011100000010101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01010011100000010101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01010011100000010110) && ({row_reg, col_reg}<20'b01010011101101110010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01010011101101110010) && ({row_reg, col_reg}<20'b01010011101101110100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01010011101101110100) && ({row_reg, col_reg}<20'b01010011101101110110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01010011101101110110) && ({row_reg, col_reg}<20'b01010011101101111000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01010011101101111000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==20'b01010011101101111001)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01010011101101111010)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01010011101101111011)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01010011101101111100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=20'b01010011101101111101) && ({row_reg, col_reg}<20'b01010011101101111111)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01010011101101111111)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01010011101110000000) && ({row_reg, col_reg}<20'b01010011110000000011)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=20'b01010011110000000011) && ({row_reg, col_reg}<20'b01010011110000000101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=20'b01010011110000000101) && ({row_reg, col_reg}<20'b01010011110000001001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01010011110000001001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=20'b01010011110000001010) && ({row_reg, col_reg}<20'b01010011110000001100)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01010011110000001100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==20'b01010011110000001101)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01010011110000001110)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==20'b01010011110000001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01010011110000010000) && ({row_reg, col_reg}<20'b01010011110000010011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01010011110000010011) && ({row_reg, col_reg}<20'b01010011110000010101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01010011110000010101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01010011110000010110) && ({row_reg, col_reg}<20'b01010011111101110011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01010011111101110011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01010011111101110100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01010011111101110101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01010011111101110110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==20'b01010011111101110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==20'b01010011111101111000)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=20'b01010011111101111001) && ({row_reg, col_reg}<20'b01010011111101111110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01010011111101111110)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01010011111101111111) && ({row_reg, col_reg}<20'b01010100000000001111)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01010100000000001111)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01010100000000010000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==20'b01010100000000010001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==20'b01010100000000010010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01010100000000010011) && ({row_reg, col_reg}<20'b01010100000000010111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01010100000000010111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01010100000000011000) && ({row_reg, col_reg}<20'b01010100000100011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01010100000100011000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01010100000100011001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01010100000100011010) && ({row_reg, col_reg}<20'b01010100000100011100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01010100000100011100) && ({row_reg, col_reg}<20'b01010100000101001010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01010100000101001010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01010100000101001011) && ({row_reg, col_reg}<20'b01010100000101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01010100000101001101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01010100000101001110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01010100000101001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01010100000101010000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01010100000101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01010100000101010010) && ({row_reg, col_reg}<20'b01010100000101010100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01010100000101010100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01010100000101010101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01010100000101010110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01010100000101010111) && ({row_reg, col_reg}<20'b01010100001000110000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01010100001000110000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01010100001000110001) && ({row_reg, col_reg}<20'b01010100001000110100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01010100001000110100) && ({row_reg, col_reg}<20'b01010100001000110110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01010100001000110110) && ({row_reg, col_reg}<20'b01010100001000111000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01010100001000111000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01010100001000111001) && ({row_reg, col_reg}<20'b01010100001000111011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01010100001000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01010100001000111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01010100001000111101) && ({row_reg, col_reg}<20'b01010100001000111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01010100001000111111) && ({row_reg, col_reg}<20'b01010100001001100001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01010100001001100001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01010100001001100010) && ({row_reg, col_reg}<20'b01010100001001101011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01010100001001101011) && ({row_reg, col_reg}<20'b01010100001001101101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01010100001001101101) && ({row_reg, col_reg}<20'b01010100001001101111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01010100001001101111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01010100001001110000) && ({row_reg, col_reg}<20'b01010100001101101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01010100001101101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01010100001101101001) && ({row_reg, col_reg}<20'b01010100001101101011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01010100001101101011) && ({row_reg, col_reg}<20'b01010100001101101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01010100001101101110) && ({row_reg, col_reg}<20'b01010100001101110100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01010100001101110100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01010100001101110101)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==20'b01010100001101110110)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==20'b01010100001101110111)) color_data = 12'b110111011101;

		if(({row_reg, col_reg}>=20'b01010100001101111000) && ({row_reg, col_reg}<20'b01010100010000001101)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01010100010000001101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=20'b01010100010000001110) && ({row_reg, col_reg}<20'b01010100010000010001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01010100010000010001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==20'b01010100010000010010)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01010100010000010011)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01010100010000010100) && ({row_reg, col_reg}<20'b01010100010000010110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=20'b01010100010000010110) && ({row_reg, col_reg}<20'b01010100010000011001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01010100010000011001) && ({row_reg, col_reg}<20'b01010100010000011101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01010100010000011101) && ({row_reg, col_reg}<20'b01010100010000011111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01010100010000011111) && ({row_reg, col_reg}<20'b01010100010100011010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01010100010100011010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01010100010100011011) && ({row_reg, col_reg}<20'b01010100010100011101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01010100010100011101) && ({row_reg, col_reg}<20'b01010100010100100000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01010100010100100000) && ({row_reg, col_reg}<20'b01010100010101001010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01010100010101001010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01010100010101001011) && ({row_reg, col_reg}<20'b01010100010101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01010100010101001101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01010100010101001110) && ({row_reg, col_reg}<20'b01010100010101010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01010100010101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01010100010101010010) && ({row_reg, col_reg}<20'b01010100010101010100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01010100010101010100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01010100010101010101) && ({row_reg, col_reg}<20'b01010100011000110010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01010100011000110010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01010100011000110011) && ({row_reg, col_reg}<20'b01010100011000110110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01010100011000110110) && ({row_reg, col_reg}<20'b01010100011000111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01010100011000111001) && ({row_reg, col_reg}<20'b01010100011000111011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01010100011000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01010100011000111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01010100011000111101) && ({row_reg, col_reg}<20'b01010100011000111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01010100011000111111) && ({row_reg, col_reg}<20'b01010100011001100001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01010100011001100001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01010100011001100010) && ({row_reg, col_reg}<20'b01010100011001100111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01010100011001100111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01010100011001101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01010100011001101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01010100011001101010) && ({row_reg, col_reg}<20'b01010100011001101110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01010100011001101110) && ({row_reg, col_reg}<20'b01010100011001110000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01010100011001110000) && ({row_reg, col_reg}<20'b01010100011101101010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01010100011101101010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01010100011101101011) && ({row_reg, col_reg}<20'b01010100011101101110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01010100011101101110) && ({row_reg, col_reg}<20'b01010100011101110000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01010100011101110000) && ({row_reg, col_reg}<20'b01010100011101110010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=20'b01010100011101110010) && ({row_reg, col_reg}<20'b01010100011101110100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==20'b01010100011101110100)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01010100011101110101)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==20'b01010100011101110110)) color_data = 12'b110111011101;

		if(({row_reg, col_reg}>=20'b01010100011101110111) && ({row_reg, col_reg}<20'b01010100100000001110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=20'b01010100100000001110) && ({row_reg, col_reg}<20'b01010100100000010001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=20'b01010100100000010001) && ({row_reg, col_reg}<20'b01010100100000010011)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01010100100000010011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01010100100000010100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=20'b01010100100000010101) && ({row_reg, col_reg}<20'b01010100100000010111)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01010100100000010111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01010100100000011000) && ({row_reg, col_reg}<20'b01010100100000011011)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=20'b01010100100000011011) && ({row_reg, col_reg}<20'b01010100100100011010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01010100100100011010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=20'b01010100100100011011) && ({row_reg, col_reg}<20'b01010100100100011101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01010100100100011101)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==20'b01010100100100011110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01010100100100011111) && ({row_reg, col_reg}<20'b01010100100101001000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01010100100101001000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01010100100101001001) && ({row_reg, col_reg}<20'b01010100100101001011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01010100100101001011) && ({row_reg, col_reg}<20'b01010100100101001101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01010100100101001101) && ({row_reg, col_reg}<20'b01010100100101001111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01010100100101001111) && ({row_reg, col_reg}<20'b01010100100101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01010100100101010001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=20'b01010100100101010010) && ({row_reg, col_reg}<20'b01010100101000110010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01010100101000110010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=20'b01010100101000110011) && ({row_reg, col_reg}<20'b01010100101000111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01010100101000111001) && ({row_reg, col_reg}<20'b01010100101000111011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01010100101000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01010100101000111100) && ({row_reg, col_reg}<20'b01010100101000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01010100101000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01010100101000111111) && ({row_reg, col_reg}<20'b01010100101001100001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01010100101001100001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01010100101001100010) && ({row_reg, col_reg}<20'b01010100101001100100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01010100101001100100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01010100101001100101) && ({row_reg, col_reg}<20'b01010100101001100111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01010100101001100111) && ({row_reg, col_reg}<20'b01010100101001101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01010100101001101001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=20'b01010100101001101010) && ({row_reg, col_reg}<20'b01010100101101101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01010100101101101100) && ({row_reg, col_reg}<20'b01010100101101101110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=20'b01010100101101101110) && ({row_reg, col_reg}<20'b01010100101101110000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==20'b01010100101101110000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01010100101101110001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==20'b01010100101101110010)) color_data = 12'b110111011101;

		if(({row_reg, col_reg}>=20'b01010100101101110011) && ({row_reg, col_reg}<20'b01010100110000010111)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=20'b01010100110000010111) && ({row_reg, col_reg}<20'b01010100110000011010)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=20'b01010100110000011010) && ({row_reg, col_reg}<20'b01010100110100011110)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==20'b01010100110100011110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==20'b01010100110100011111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01010100110100100000) && ({row_reg, col_reg}<20'b01010100110101001000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01010100110101001000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01010100110101001001) && ({row_reg, col_reg}<20'b01010100110101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01010100110101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01010100110101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01010100110101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01010100110101001111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=20'b01010100110101010000) && ({row_reg, col_reg}<20'b01010100111000110110)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==20'b01010100111000110110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01010100111000110111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==20'b01010100111000111000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01010100111000111001) && ({row_reg, col_reg}<20'b01010100111000111011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01010100111000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01010100111000111100) && ({row_reg, col_reg}<20'b01010100111000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01010100111000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01010100111000111111) && ({row_reg, col_reg}<20'b01010100111001100100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01010100111001100100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01010100111001100101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01010100111001100110) && ({row_reg, col_reg}<20'b01010100111001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01010100111001101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01010100111001101001) && ({row_reg, col_reg}<20'b01010100111101101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=20'b01010100111101101100) && ({row_reg, col_reg}<20'b01010100111101101110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=20'b01010100111101101110) && ({row_reg, col_reg}<20'b01010100111101110101)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01010100111101110101)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01010100111101110110) && ({row_reg, col_reg}<20'b01010101000000001011)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01010101000000001011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=20'b01010101000000001100) && ({row_reg, col_reg}<20'b01010101000000010111)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=20'b01010101000000010111) && ({row_reg, col_reg}<20'b01010101000000011001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=20'b01010101000000011001) && ({row_reg, col_reg}<20'b01010101000100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01010101000100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01010101000100011111) && ({row_reg, col_reg}<20'b01010101000101001000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01010101000101001000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01010101000101001001) && ({row_reg, col_reg}<20'b01010101000101001110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01010101000101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01010101000101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==20'b01010101000101010000)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=20'b01010101000101010001) && ({row_reg, col_reg}<20'b01010101001000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01010101001000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01010101001000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01010101001000111000) && ({row_reg, col_reg}<20'b01010101001000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01010101001000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01010101001000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01010101001000111100) && ({row_reg, col_reg}<20'b01010101001001100100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01010101001001100100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01010101001001100101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01010101001001100110) && ({row_reg, col_reg}<20'b01010101001001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01010101001001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01010101001001101001) && ({row_reg, col_reg}<20'b01010101001101101101)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01010101001101101101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=20'b01010101001101101110) && ({row_reg, col_reg}<20'b01010101001101110000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01010101001101110000)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01010101001101110001) && ({row_reg, col_reg}<20'b01010101010100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01010101010100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01010101010100011111) && ({row_reg, col_reg}<20'b01010101010101001010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01010101010101001010) && ({row_reg, col_reg}<20'b01010101010101001101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01010101010101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01010101010101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01010101010101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01010101010101010000) && ({row_reg, col_reg}<20'b01010101011000110011)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01010101011000110011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=20'b01010101011000110100) && ({row_reg, col_reg}<20'b01010101011000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01010101011000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01010101011000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01010101011000111000) && ({row_reg, col_reg}<20'b01010101011000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01010101011000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01010101011000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01010101011000111100) && ({row_reg, col_reg}<20'b01010101011001100100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01010101011001100100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01010101011001100101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01010101011001100110) && ({row_reg, col_reg}<20'b01010101011001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01010101011001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01010101011001101001) && ({row_reg, col_reg}<20'b01010101011101110010)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=20'b01010101011101110010) && ({row_reg, col_reg}<20'b01010101011101110101)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01010101011101110101) && ({row_reg, col_reg}<20'b01010101100100011001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01010101100100011001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=20'b01010101100100011010) && ({row_reg, col_reg}<20'b01010101100100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01010101100100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01010101100100011111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01010101100100100000) && ({row_reg, col_reg}<20'b01010101100101001001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01010101100101001001) && ({row_reg, col_reg}<20'b01010101100101001011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01010101100101001011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01010101100101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01010101100101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01010101100101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01010101100101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01010101100101010000) && ({row_reg, col_reg}<20'b01010101100101010110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01010101100101010110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=20'b01010101100101010111) && ({row_reg, col_reg}<20'b01010101101000110011)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01010101101000110011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==20'b01010101101000110100)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01010101101000110101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==20'b01010101101000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01010101101000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01010101101000111000) && ({row_reg, col_reg}<20'b01010101101000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01010101101000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01010101101000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01010101101000111100) && ({row_reg, col_reg}<20'b01010101101000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01010101101000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01010101101000111111) && ({row_reg, col_reg}<20'b01010101101001100100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01010101101001100100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01010101101001100101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01010101101001100110) && ({row_reg, col_reg}<20'b01010101101001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01010101101001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01010101101001101001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=20'b01010101101001101010) && ({row_reg, col_reg}<20'b01010101101001101111)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01010101101001101111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=20'b01010101101001110000) && ({row_reg, col_reg}<20'b01010101101101101010)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01010101101101101010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=20'b01010101101101101011) && ({row_reg, col_reg}<20'b01010101101101101111)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=20'b01010101101101101111) && ({row_reg, col_reg}<20'b01010101101101110001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=20'b01010101101101110001) && ({row_reg, col_reg}<20'b01010101101101110111)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01010101101101110111)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01010101101101111000) && ({row_reg, col_reg}<20'b01010101110000001101)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01010101110000001101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=20'b01010101110000001110) && ({row_reg, col_reg}<20'b01010101110100011001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01010101110100011001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=20'b01010101110100011010) && ({row_reg, col_reg}<20'b01010101110100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01010101110100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01010101110100011111) && ({row_reg, col_reg}<20'b01010101110101001001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01010101110101001001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01010101110101001010) && ({row_reg, col_reg}<20'b01010101110101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01010101110101001100) && ({row_reg, col_reg}<20'b01010101110101001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01010101110101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01010101110101010000) && ({row_reg, col_reg}<20'b01010101111000110000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01010101111000110000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=20'b01010101111000110001) && ({row_reg, col_reg}<20'b01010101111000110011)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01010101111000110011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==20'b01010101111000110100)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01010101111000110101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==20'b01010101111000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01010101111000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==20'b01010101111000111000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01010101111000111001) && ({row_reg, col_reg}<20'b01010101111000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01010101111000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01010101111000111111) && ({row_reg, col_reg}<20'b01010101111001100100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01010101111001100100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01010101111001100101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01010101111001100110) && ({row_reg, col_reg}<20'b01010101111001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01010101111001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01010101111001101001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=20'b01010101111001101010) && ({row_reg, col_reg}<20'b01010101111001101101)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01010101111001101101)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01010101111001101110) && ({row_reg, col_reg}<20'b01010110000100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01010110000100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01010110000100011111) && ({row_reg, col_reg}<20'b01010110000101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01010110000101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01010110000101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01010110000101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01010110000101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01010110000101010000) && ({row_reg, col_reg}<20'b01010110001000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01010110001000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01010110001000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01010110001000111000) && ({row_reg, col_reg}<20'b01010110001000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01010110001000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01010110001000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01010110001000111100) && ({row_reg, col_reg}<20'b01010110001000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01010110001000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01010110001000111111) && ({row_reg, col_reg}<20'b01010110001001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01010110001001100110) && ({row_reg, col_reg}<20'b01010110001001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01010110001001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01010110001001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01010110001001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01010110001001101011) && ({row_reg, col_reg}<20'b01010110010100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01010110010100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01010110010100011111) && ({row_reg, col_reg}<20'b01010110010101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01010110010101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01010110010101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01010110010101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01010110010101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01010110010101010000) && ({row_reg, col_reg}<20'b01010110011000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01010110011000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01010110011000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01010110011000111000) && ({row_reg, col_reg}<20'b01010110011000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01010110011000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01010110011000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01010110011000111100) && ({row_reg, col_reg}<20'b01010110011000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01010110011000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01010110011000111111) && ({row_reg, col_reg}<20'b01010110011001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01010110011001100110) && ({row_reg, col_reg}<20'b01010110011001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01010110011001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01010110011001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01010110011001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01010110011001101011) && ({row_reg, col_reg}<20'b01010110100100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01010110100100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01010110100100011111) && ({row_reg, col_reg}<20'b01010110100101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01010110100101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01010110100101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01010110100101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01010110100101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01010110100101010000) && ({row_reg, col_reg}<20'b01010110101000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01010110101000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01010110101000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01010110101000111000) && ({row_reg, col_reg}<20'b01010110101000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01010110101000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01010110101000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01010110101000111100) && ({row_reg, col_reg}<20'b01010110101000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01010110101000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01010110101000111111) && ({row_reg, col_reg}<20'b01010110101001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01010110101001100110) && ({row_reg, col_reg}<20'b01010110101001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01010110101001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01010110101001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01010110101001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01010110101001101011) && ({row_reg, col_reg}<20'b01010110110100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01010110110100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01010110110100011111) && ({row_reg, col_reg}<20'b01010110110101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01010110110101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01010110110101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01010110110101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01010110110101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01010110110101010000) && ({row_reg, col_reg}<20'b01010110111000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01010110111000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01010110111000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01010110111000111000) && ({row_reg, col_reg}<20'b01010110111000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01010110111000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01010110111000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01010110111000111100) && ({row_reg, col_reg}<20'b01010110111000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01010110111000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01010110111000111111) && ({row_reg, col_reg}<20'b01010110111001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01010110111001100110) && ({row_reg, col_reg}<20'b01010110111001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01010110111001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01010110111001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01010110111001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01010110111001101011) && ({row_reg, col_reg}<20'b01010111000100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01010111000100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01010111000100011111) && ({row_reg, col_reg}<20'b01010111000101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01010111000101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01010111000101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01010111000101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01010111000101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01010111000101010000) && ({row_reg, col_reg}<20'b01010111001000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01010111001000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01010111001000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01010111001000111000) && ({row_reg, col_reg}<20'b01010111001000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01010111001000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01010111001000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01010111001000111100) && ({row_reg, col_reg}<20'b01010111001000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01010111001000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01010111001000111111) && ({row_reg, col_reg}<20'b01010111001001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01010111001001100110) && ({row_reg, col_reg}<20'b01010111001001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01010111001001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01010111001001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01010111001001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01010111001001101011) && ({row_reg, col_reg}<20'b01010111010100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01010111010100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01010111010100011111) && ({row_reg, col_reg}<20'b01010111010101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01010111010101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01010111010101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01010111010101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01010111010101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01010111010101010000) && ({row_reg, col_reg}<20'b01010111011000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01010111011000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01010111011000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01010111011000111000) && ({row_reg, col_reg}<20'b01010111011000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01010111011000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01010111011000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01010111011000111100) && ({row_reg, col_reg}<20'b01010111011000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01010111011000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01010111011000111111) && ({row_reg, col_reg}<20'b01010111011001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01010111011001100110) && ({row_reg, col_reg}<20'b01010111011001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01010111011001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01010111011001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01010111011001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01010111011001101011) && ({row_reg, col_reg}<20'b01010111100100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01010111100100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01010111100100011111) && ({row_reg, col_reg}<20'b01010111100101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01010111100101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01010111100101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01010111100101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01010111100101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01010111100101010000) && ({row_reg, col_reg}<20'b01010111101000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01010111101000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01010111101000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01010111101000111000) && ({row_reg, col_reg}<20'b01010111101000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01010111101000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01010111101000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01010111101000111100) && ({row_reg, col_reg}<20'b01010111101000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01010111101000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01010111101000111111) && ({row_reg, col_reg}<20'b01010111101001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01010111101001100110) && ({row_reg, col_reg}<20'b01010111101001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01010111101001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01010111101001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01010111101001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01010111101001101011) && ({row_reg, col_reg}<20'b01010111110100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01010111110100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01010111110100011111) && ({row_reg, col_reg}<20'b01010111110101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01010111110101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01010111110101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01010111110101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01010111110101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01010111110101010000) && ({row_reg, col_reg}<20'b01010111111000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01010111111000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01010111111000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01010111111000111000) && ({row_reg, col_reg}<20'b01010111111000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01010111111000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01010111111000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01010111111000111100) && ({row_reg, col_reg}<20'b01010111111000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01010111111000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01010111111000111111) && ({row_reg, col_reg}<20'b01010111111001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01010111111001100110) && ({row_reg, col_reg}<20'b01010111111001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01010111111001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01010111111001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01010111111001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01010111111001101011) && ({row_reg, col_reg}<20'b01011000000100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01011000000100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01011000000100011111) && ({row_reg, col_reg}<20'b01011000000101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01011000000101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01011000000101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01011000000101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01011000000101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01011000000101010000) && ({row_reg, col_reg}<20'b01011000001000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01011000001000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01011000001000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01011000001000111000) && ({row_reg, col_reg}<20'b01011000001000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01011000001000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01011000001000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01011000001000111100) && ({row_reg, col_reg}<20'b01011000001000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01011000001000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01011000001000111111) && ({row_reg, col_reg}<20'b01011000001001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01011000001001100110) && ({row_reg, col_reg}<20'b01011000001001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01011000001001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01011000001001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01011000001001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01011000001001101011) && ({row_reg, col_reg}<20'b01011000010100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01011000010100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01011000010100011111) && ({row_reg, col_reg}<20'b01011000010101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01011000010101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01011000010101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01011000010101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01011000010101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01011000010101010000) && ({row_reg, col_reg}<20'b01011000011000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01011000011000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01011000011000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01011000011000111000) && ({row_reg, col_reg}<20'b01011000011000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01011000011000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01011000011000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01011000011000111100) && ({row_reg, col_reg}<20'b01011000011000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01011000011000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01011000011000111111) && ({row_reg, col_reg}<20'b01011000011001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01011000011001100110) && ({row_reg, col_reg}<20'b01011000011001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01011000011001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01011000011001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01011000011001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01011000011001101011) && ({row_reg, col_reg}<20'b01011000100100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01011000100100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01011000100100011111) && ({row_reg, col_reg}<20'b01011000100101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01011000100101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01011000100101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01011000100101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01011000100101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01011000100101010000) && ({row_reg, col_reg}<20'b01011000101000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01011000101000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01011000101000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01011000101000111000) && ({row_reg, col_reg}<20'b01011000101000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01011000101000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01011000101000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01011000101000111100) && ({row_reg, col_reg}<20'b01011000101000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01011000101000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01011000101000111111) && ({row_reg, col_reg}<20'b01011000101001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01011000101001100110) && ({row_reg, col_reg}<20'b01011000101001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01011000101001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01011000101001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01011000101001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01011000101001101011) && ({row_reg, col_reg}<20'b01011000110100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01011000110100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01011000110100011111) && ({row_reg, col_reg}<20'b01011000110101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01011000110101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01011000110101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01011000110101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01011000110101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01011000110101010000) && ({row_reg, col_reg}<20'b01011000111000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01011000111000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01011000111000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01011000111000111000) && ({row_reg, col_reg}<20'b01011000111000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01011000111000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01011000111000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01011000111000111100) && ({row_reg, col_reg}<20'b01011000111000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01011000111000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01011000111000111111) && ({row_reg, col_reg}<20'b01011000111001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01011000111001100110) && ({row_reg, col_reg}<20'b01011000111001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01011000111001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01011000111001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01011000111001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01011000111001101011) && ({row_reg, col_reg}<20'b01011001000100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01011001000100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01011001000100011111) && ({row_reg, col_reg}<20'b01011001000101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01011001000101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01011001000101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01011001000101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01011001000101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01011001000101010000) && ({row_reg, col_reg}<20'b01011001001000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01011001001000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01011001001000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01011001001000111000) && ({row_reg, col_reg}<20'b01011001001000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01011001001000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01011001001000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01011001001000111100) && ({row_reg, col_reg}<20'b01011001001000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01011001001000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01011001001000111111) && ({row_reg, col_reg}<20'b01011001001001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01011001001001100110) && ({row_reg, col_reg}<20'b01011001001001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01011001001001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01011001001001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01011001001001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01011001001001101011) && ({row_reg, col_reg}<20'b01011001010100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01011001010100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01011001010100011111) && ({row_reg, col_reg}<20'b01011001010101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01011001010101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01011001010101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01011001010101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01011001010101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01011001010101010000) && ({row_reg, col_reg}<20'b01011001011000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01011001011000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01011001011000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01011001011000111000) && ({row_reg, col_reg}<20'b01011001011000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01011001011000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01011001011000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01011001011000111100) && ({row_reg, col_reg}<20'b01011001011000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01011001011000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01011001011000111111) && ({row_reg, col_reg}<20'b01011001011001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01011001011001100110) && ({row_reg, col_reg}<20'b01011001011001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01011001011001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01011001011001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01011001011001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01011001011001101011) && ({row_reg, col_reg}<20'b01011001100100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01011001100100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01011001100100011111) && ({row_reg, col_reg}<20'b01011001100101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01011001100101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01011001100101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01011001100101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01011001100101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01011001100101010000) && ({row_reg, col_reg}<20'b01011001101000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01011001101000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01011001101000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01011001101000111000) && ({row_reg, col_reg}<20'b01011001101000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01011001101000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01011001101000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01011001101000111100) && ({row_reg, col_reg}<20'b01011001101000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01011001101000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01011001101000111111) && ({row_reg, col_reg}<20'b01011001101001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01011001101001100110) && ({row_reg, col_reg}<20'b01011001101001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01011001101001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01011001101001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01011001101001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01011001101001101011) && ({row_reg, col_reg}<20'b01011001110100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01011001110100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01011001110100011111) && ({row_reg, col_reg}<20'b01011001110101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01011001110101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01011001110101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01011001110101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01011001110101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01011001110101010000) && ({row_reg, col_reg}<20'b01011001111000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01011001111000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01011001111000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01011001111000111000) && ({row_reg, col_reg}<20'b01011001111000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01011001111000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01011001111000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01011001111000111100) && ({row_reg, col_reg}<20'b01011001111000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01011001111000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01011001111000111111) && ({row_reg, col_reg}<20'b01011001111001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01011001111001100110) && ({row_reg, col_reg}<20'b01011001111001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01011001111001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01011001111001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01011001111001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01011001111001101011) && ({row_reg, col_reg}<20'b01011010000100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01011010000100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01011010000100011111) && ({row_reg, col_reg}<20'b01011010000101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01011010000101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01011010000101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01011010000101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01011010000101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01011010000101010000) && ({row_reg, col_reg}<20'b01011010001000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01011010001000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01011010001000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01011010001000111000) && ({row_reg, col_reg}<20'b01011010001000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01011010001000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01011010001000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01011010001000111100) && ({row_reg, col_reg}<20'b01011010001000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01011010001000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01011010001000111111) && ({row_reg, col_reg}<20'b01011010001001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01011010001001100110) && ({row_reg, col_reg}<20'b01011010001001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01011010001001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01011010001001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01011010001001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01011010001001101011) && ({row_reg, col_reg}<20'b01011010010100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01011010010100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01011010010100011111) && ({row_reg, col_reg}<20'b01011010010101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01011010010101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01011010010101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01011010010101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01011010010101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01011010010101010000) && ({row_reg, col_reg}<20'b01011010011000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01011010011000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01011010011000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01011010011000111000) && ({row_reg, col_reg}<20'b01011010011000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01011010011000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01011010011000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01011010011000111100) && ({row_reg, col_reg}<20'b01011010011000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01011010011000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01011010011000111111) && ({row_reg, col_reg}<20'b01011010011001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01011010011001100110) && ({row_reg, col_reg}<20'b01011010011001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01011010011001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01011010011001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01011010011001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01011010011001101011) && ({row_reg, col_reg}<20'b01011010100100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01011010100100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01011010100100011111) && ({row_reg, col_reg}<20'b01011010100101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01011010100101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01011010100101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01011010100101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01011010100101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01011010100101010000) && ({row_reg, col_reg}<20'b01011010101000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01011010101000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01011010101000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01011010101000111000) && ({row_reg, col_reg}<20'b01011010101000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01011010101000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01011010101000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01011010101000111100) && ({row_reg, col_reg}<20'b01011010101000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01011010101000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01011010101000111111) && ({row_reg, col_reg}<20'b01011010101001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01011010101001100110) && ({row_reg, col_reg}<20'b01011010101001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01011010101001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01011010101001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01011010101001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01011010101001101011) && ({row_reg, col_reg}<20'b01011010110100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01011010110100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01011010110100011111) && ({row_reg, col_reg}<20'b01011010110101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01011010110101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01011010110101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01011010110101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01011010110101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01011010110101010000) && ({row_reg, col_reg}<20'b01011010111000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01011010111000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01011010111000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01011010111000111000) && ({row_reg, col_reg}<20'b01011010111000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01011010111000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01011010111000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01011010111000111100) && ({row_reg, col_reg}<20'b01011010111000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01011010111000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01011010111000111111) && ({row_reg, col_reg}<20'b01011010111001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01011010111001100110) && ({row_reg, col_reg}<20'b01011010111001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01011010111001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01011010111001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01011010111001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01011010111001101011) && ({row_reg, col_reg}<20'b01011011000100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01011011000100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01011011000100011111) && ({row_reg, col_reg}<20'b01011011000101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01011011000101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01011011000101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01011011000101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01011011000101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01011011000101010000) && ({row_reg, col_reg}<20'b01011011001000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01011011001000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01011011001000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01011011001000111000) && ({row_reg, col_reg}<20'b01011011001000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01011011001000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01011011001000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01011011001000111100) && ({row_reg, col_reg}<20'b01011011001000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01011011001000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01011011001000111111) && ({row_reg, col_reg}<20'b01011011001001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01011011001001100110) && ({row_reg, col_reg}<20'b01011011001001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01011011001001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01011011001001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01011011001001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01011011001001101011) && ({row_reg, col_reg}<20'b01011011010100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01011011010100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01011011010100011111) && ({row_reg, col_reg}<20'b01011011010101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01011011010101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01011011010101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01011011010101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01011011010101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01011011010101010000) && ({row_reg, col_reg}<20'b01011011011000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01011011011000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01011011011000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01011011011000111000) && ({row_reg, col_reg}<20'b01011011011000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01011011011000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01011011011000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01011011011000111100) && ({row_reg, col_reg}<20'b01011011011000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01011011011000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01011011011000111111) && ({row_reg, col_reg}<20'b01011011011001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01011011011001100110) && ({row_reg, col_reg}<20'b01011011011001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01011011011001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01011011011001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01011011011001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01011011011001101011) && ({row_reg, col_reg}<20'b01011011100100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01011011100100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01011011100100011111) && ({row_reg, col_reg}<20'b01011011100101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01011011100101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01011011100101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01011011100101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01011011100101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01011011100101010000) && ({row_reg, col_reg}<20'b01011011101000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01011011101000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01011011101000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01011011101000111000) && ({row_reg, col_reg}<20'b01011011101000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01011011101000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01011011101000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01011011101000111100) && ({row_reg, col_reg}<20'b01011011101000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01011011101000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01011011101000111111) && ({row_reg, col_reg}<20'b01011011101001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01011011101001100110) && ({row_reg, col_reg}<20'b01011011101001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01011011101001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01011011101001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01011011101001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01011011101001101011) && ({row_reg, col_reg}<20'b01011011110100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01011011110100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01011011110100011111) && ({row_reg, col_reg}<20'b01011011110101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01011011110101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01011011110101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01011011110101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01011011110101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01011011110101010000) && ({row_reg, col_reg}<20'b01011011111000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01011011111000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01011011111000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01011011111000111000) && ({row_reg, col_reg}<20'b01011011111000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01011011111000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01011011111000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01011011111000111100) && ({row_reg, col_reg}<20'b01011011111000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01011011111000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01011011111000111111) && ({row_reg, col_reg}<20'b01011011111001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01011011111001100110) && ({row_reg, col_reg}<20'b01011011111001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01011011111001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01011011111001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01011011111001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01011011111001101011) && ({row_reg, col_reg}<20'b01011100000100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01011100000100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01011100000100011111) && ({row_reg, col_reg}<20'b01011100000101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01011100000101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01011100000101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01011100000101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01011100000101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01011100000101010000) && ({row_reg, col_reg}<20'b01011100001000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01011100001000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01011100001000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01011100001000111000) && ({row_reg, col_reg}<20'b01011100001000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01011100001000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01011100001000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01011100001000111100) && ({row_reg, col_reg}<20'b01011100001000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01011100001000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01011100001000111111) && ({row_reg, col_reg}<20'b01011100001001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01011100001001100110) && ({row_reg, col_reg}<20'b01011100001001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01011100001001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01011100001001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01011100001001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01011100001001101011) && ({row_reg, col_reg}<20'b01011100010100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01011100010100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01011100010100011111) && ({row_reg, col_reg}<20'b01011100010101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01011100010101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01011100010101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01011100010101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01011100010101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01011100010101010000) && ({row_reg, col_reg}<20'b01011100011000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01011100011000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01011100011000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01011100011000111000) && ({row_reg, col_reg}<20'b01011100011000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01011100011000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01011100011000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01011100011000111100) && ({row_reg, col_reg}<20'b01011100011000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01011100011000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01011100011000111111) && ({row_reg, col_reg}<20'b01011100011001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01011100011001100110) && ({row_reg, col_reg}<20'b01011100011001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01011100011001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01011100011001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01011100011001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01011100011001101011) && ({row_reg, col_reg}<20'b01011100100100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01011100100100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01011100100100011111) && ({row_reg, col_reg}<20'b01011100100101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01011100100101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01011100100101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01011100100101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01011100100101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01011100100101010000) && ({row_reg, col_reg}<20'b01011100101000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01011100101000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01011100101000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01011100101000111000) && ({row_reg, col_reg}<20'b01011100101000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01011100101000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01011100101000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01011100101000111100) && ({row_reg, col_reg}<20'b01011100101000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01011100101000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01011100101000111111) && ({row_reg, col_reg}<20'b01011100101001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01011100101001100110) && ({row_reg, col_reg}<20'b01011100101001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01011100101001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01011100101001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01011100101001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01011100101001101011) && ({row_reg, col_reg}<20'b01011100110100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01011100110100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01011100110100011111) && ({row_reg, col_reg}<20'b01011100110101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01011100110101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01011100110101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01011100110101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01011100110101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01011100110101010000) && ({row_reg, col_reg}<20'b01011100111000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01011100111000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01011100111000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01011100111000111000) && ({row_reg, col_reg}<20'b01011100111000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01011100111000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01011100111000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01011100111000111100) && ({row_reg, col_reg}<20'b01011100111000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01011100111000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01011100111000111111) && ({row_reg, col_reg}<20'b01011100111001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01011100111001100110) && ({row_reg, col_reg}<20'b01011100111001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01011100111001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01011100111001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01011100111001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01011100111001101011) && ({row_reg, col_reg}<20'b01011101000100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01011101000100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01011101000100011111) && ({row_reg, col_reg}<20'b01011101000101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01011101000101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01011101000101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01011101000101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01011101000101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01011101000101010000) && ({row_reg, col_reg}<20'b01011101001000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01011101001000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01011101001000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01011101001000111000) && ({row_reg, col_reg}<20'b01011101001000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01011101001000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01011101001000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01011101001000111100) && ({row_reg, col_reg}<20'b01011101001000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01011101001000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01011101001000111111) && ({row_reg, col_reg}<20'b01011101001001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01011101001001100110) && ({row_reg, col_reg}<20'b01011101001001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01011101001001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01011101001001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01011101001001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01011101001001101011) && ({row_reg, col_reg}<20'b01011101010100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01011101010100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01011101010100011111) && ({row_reg, col_reg}<20'b01011101010101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01011101010101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01011101010101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01011101010101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01011101010101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01011101010101010000) && ({row_reg, col_reg}<20'b01011101011000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01011101011000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01011101011000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01011101011000111000) && ({row_reg, col_reg}<20'b01011101011000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01011101011000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01011101011000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01011101011000111100) && ({row_reg, col_reg}<20'b01011101011000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01011101011000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01011101011000111111) && ({row_reg, col_reg}<20'b01011101011001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01011101011001100110) && ({row_reg, col_reg}<20'b01011101011001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01011101011001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01011101011001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01011101011001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01011101011001101011) && ({row_reg, col_reg}<20'b01011101100100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01011101100100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01011101100100011111) && ({row_reg, col_reg}<20'b01011101100101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01011101100101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01011101100101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01011101100101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01011101100101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01011101100101010000) && ({row_reg, col_reg}<20'b01011101101000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01011101101000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01011101101000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01011101101000111000) && ({row_reg, col_reg}<20'b01011101101000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01011101101000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01011101101000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01011101101000111100) && ({row_reg, col_reg}<20'b01011101101000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01011101101000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01011101101000111111) && ({row_reg, col_reg}<20'b01011101101001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01011101101001100110) && ({row_reg, col_reg}<20'b01011101101001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01011101101001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01011101101001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01011101101001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01011101101001101011) && ({row_reg, col_reg}<20'b01011101110100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01011101110100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01011101110100011111) && ({row_reg, col_reg}<20'b01011101110101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01011101110101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01011101110101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01011101110101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01011101110101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01011101110101010000) && ({row_reg, col_reg}<20'b01011101111000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01011101111000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01011101111000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01011101111000111000) && ({row_reg, col_reg}<20'b01011101111000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01011101111000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01011101111000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01011101111000111100) && ({row_reg, col_reg}<20'b01011101111000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01011101111000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01011101111000111111) && ({row_reg, col_reg}<20'b01011101111001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01011101111001100110) && ({row_reg, col_reg}<20'b01011101111001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01011101111001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01011101111001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01011101111001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01011101111001101011) && ({row_reg, col_reg}<20'b01011110000100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01011110000100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01011110000100011111) && ({row_reg, col_reg}<20'b01011110000101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01011110000101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01011110000101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01011110000101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01011110000101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01011110000101010000) && ({row_reg, col_reg}<20'b01011110001000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01011110001000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01011110001000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01011110001000111000) && ({row_reg, col_reg}<20'b01011110001000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01011110001000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01011110001000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01011110001000111100) && ({row_reg, col_reg}<20'b01011110001000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01011110001000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01011110001000111111) && ({row_reg, col_reg}<20'b01011110001001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01011110001001100110) && ({row_reg, col_reg}<20'b01011110001001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01011110001001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01011110001001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01011110001001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01011110001001101011) && ({row_reg, col_reg}<20'b01011110010100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01011110010100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01011110010100011111) && ({row_reg, col_reg}<20'b01011110010101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01011110010101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01011110010101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01011110010101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01011110010101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01011110010101010000) && ({row_reg, col_reg}<20'b01011110011000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01011110011000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01011110011000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01011110011000111000) && ({row_reg, col_reg}<20'b01011110011000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01011110011000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01011110011000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01011110011000111100) && ({row_reg, col_reg}<20'b01011110011000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01011110011000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01011110011000111111) && ({row_reg, col_reg}<20'b01011110011001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01011110011001100110) && ({row_reg, col_reg}<20'b01011110011001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01011110011001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01011110011001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01011110011001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01011110011001101011) && ({row_reg, col_reg}<20'b01011110100100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01011110100100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01011110100100011111) && ({row_reg, col_reg}<20'b01011110100101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01011110100101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01011110100101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01011110100101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01011110100101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01011110100101010000) && ({row_reg, col_reg}<20'b01011110101000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01011110101000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01011110101000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01011110101000111000) && ({row_reg, col_reg}<20'b01011110101000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01011110101000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01011110101000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01011110101000111100) && ({row_reg, col_reg}<20'b01011110101000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01011110101000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01011110101000111111) && ({row_reg, col_reg}<20'b01011110101001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01011110101001100110) && ({row_reg, col_reg}<20'b01011110101001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01011110101001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01011110101001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01011110101001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01011110101001101011) && ({row_reg, col_reg}<20'b01011110110100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01011110110100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01011110110100011111) && ({row_reg, col_reg}<20'b01011110110101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01011110110101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01011110110101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01011110110101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01011110110101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01011110110101010000) && ({row_reg, col_reg}<20'b01011110111000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01011110111000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01011110111000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01011110111000111000) && ({row_reg, col_reg}<20'b01011110111000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01011110111000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01011110111000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01011110111000111100) && ({row_reg, col_reg}<20'b01011110111000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01011110111000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01011110111000111111) && ({row_reg, col_reg}<20'b01011110111001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01011110111001100110) && ({row_reg, col_reg}<20'b01011110111001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01011110111001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01011110111001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01011110111001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01011110111001101011) && ({row_reg, col_reg}<20'b01011111000100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01011111000100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01011111000100011111) && ({row_reg, col_reg}<20'b01011111000101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01011111000101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01011111000101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01011111000101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01011111000101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01011111000101010000) && ({row_reg, col_reg}<20'b01011111001000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01011111001000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01011111001000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01011111001000111000) && ({row_reg, col_reg}<20'b01011111001000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01011111001000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01011111001000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01011111001000111100) && ({row_reg, col_reg}<20'b01011111001000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01011111001000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01011111001000111111) && ({row_reg, col_reg}<20'b01011111001001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01011111001001100110) && ({row_reg, col_reg}<20'b01011111001001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01011111001001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01011111001001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01011111001001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01011111001001101011) && ({row_reg, col_reg}<20'b01011111010100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01011111010100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01011111010100011111) && ({row_reg, col_reg}<20'b01011111010101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01011111010101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01011111010101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01011111010101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01011111010101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01011111010101010000) && ({row_reg, col_reg}<20'b01011111011000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01011111011000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01011111011000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01011111011000111000) && ({row_reg, col_reg}<20'b01011111011000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01011111011000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01011111011000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01011111011000111100) && ({row_reg, col_reg}<20'b01011111011000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01011111011000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01011111011000111111) && ({row_reg, col_reg}<20'b01011111011001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01011111011001100110) && ({row_reg, col_reg}<20'b01011111011001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01011111011001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01011111011001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01011111011001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01011111011001101011) && ({row_reg, col_reg}<20'b01011111100100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01011111100100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01011111100100011111) && ({row_reg, col_reg}<20'b01011111100101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01011111100101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01011111100101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01011111100101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01011111100101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01011111100101010000) && ({row_reg, col_reg}<20'b01011111101000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01011111101000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01011111101000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01011111101000111000) && ({row_reg, col_reg}<20'b01011111101000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01011111101000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01011111101000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01011111101000111100) && ({row_reg, col_reg}<20'b01011111101000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01011111101000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01011111101000111111) && ({row_reg, col_reg}<20'b01011111101001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01011111101001100110) && ({row_reg, col_reg}<20'b01011111101001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01011111101001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01011111101001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01011111101001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01011111101001101011) && ({row_reg, col_reg}<20'b01011111110100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01011111110100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01011111110100011111) && ({row_reg, col_reg}<20'b01011111110101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01011111110101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01011111110101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01011111110101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01011111110101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01011111110101010000) && ({row_reg, col_reg}<20'b01011111111000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01011111111000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01011111111000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01011111111000111000) && ({row_reg, col_reg}<20'b01011111111000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01011111111000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01011111111000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01011111111000111100) && ({row_reg, col_reg}<20'b01011111111000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01011111111000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01011111111000111111) && ({row_reg, col_reg}<20'b01011111111001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01011111111001100110) && ({row_reg, col_reg}<20'b01011111111001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01011111111001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01011111111001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01011111111001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01011111111001101011) && ({row_reg, col_reg}<20'b01100000000100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01100000000100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01100000000100011111) && ({row_reg, col_reg}<20'b01100000000101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01100000000101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01100000000101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01100000000101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01100000000101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01100000000101010000) && ({row_reg, col_reg}<20'b01100000001000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01100000001000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01100000001000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01100000001000111000) && ({row_reg, col_reg}<20'b01100000001000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01100000001000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01100000001000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01100000001000111100) && ({row_reg, col_reg}<20'b01100000001000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01100000001000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01100000001000111111) && ({row_reg, col_reg}<20'b01100000001001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01100000001001100110) && ({row_reg, col_reg}<20'b01100000001001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01100000001001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01100000001001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01100000001001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01100000001001101011) && ({row_reg, col_reg}<20'b01100000010100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01100000010100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01100000010100011111) && ({row_reg, col_reg}<20'b01100000010101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01100000010101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01100000010101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01100000010101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01100000010101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01100000010101010000) && ({row_reg, col_reg}<20'b01100000011000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01100000011000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01100000011000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01100000011000111000) && ({row_reg, col_reg}<20'b01100000011000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01100000011000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01100000011000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01100000011000111100) && ({row_reg, col_reg}<20'b01100000011000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01100000011000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01100000011000111111) && ({row_reg, col_reg}<20'b01100000011001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01100000011001100110) && ({row_reg, col_reg}<20'b01100000011001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01100000011001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01100000011001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01100000011001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01100000011001101011) && ({row_reg, col_reg}<20'b01100000100100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01100000100100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01100000100100011111) && ({row_reg, col_reg}<20'b01100000100101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01100000100101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01100000100101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01100000100101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01100000100101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01100000100101010000) && ({row_reg, col_reg}<20'b01100000101000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01100000101000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01100000101000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01100000101000111000) && ({row_reg, col_reg}<20'b01100000101000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01100000101000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01100000101000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01100000101000111100) && ({row_reg, col_reg}<20'b01100000101000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01100000101000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01100000101000111111) && ({row_reg, col_reg}<20'b01100000101001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01100000101001100110) && ({row_reg, col_reg}<20'b01100000101001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01100000101001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01100000101001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01100000101001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01100000101001101011) && ({row_reg, col_reg}<20'b01100000110100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01100000110100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01100000110100011111) && ({row_reg, col_reg}<20'b01100000110101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01100000110101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01100000110101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01100000110101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01100000110101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01100000110101010000) && ({row_reg, col_reg}<20'b01100000111000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01100000111000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01100000111000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01100000111000111000) && ({row_reg, col_reg}<20'b01100000111000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01100000111000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01100000111000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01100000111000111100) && ({row_reg, col_reg}<20'b01100000111000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01100000111000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01100000111000111111) && ({row_reg, col_reg}<20'b01100000111001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01100000111001100110) && ({row_reg, col_reg}<20'b01100000111001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01100000111001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01100000111001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01100000111001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01100000111001101011) && ({row_reg, col_reg}<20'b01100001000100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01100001000100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01100001000100011111) && ({row_reg, col_reg}<20'b01100001000101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01100001000101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01100001000101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01100001000101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01100001000101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01100001000101010000) && ({row_reg, col_reg}<20'b01100001001000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01100001001000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01100001001000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01100001001000111000) && ({row_reg, col_reg}<20'b01100001001000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01100001001000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01100001001000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01100001001000111100) && ({row_reg, col_reg}<20'b01100001001000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01100001001000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01100001001000111111) && ({row_reg, col_reg}<20'b01100001001001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01100001001001100110) && ({row_reg, col_reg}<20'b01100001001001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01100001001001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01100001001001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01100001001001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01100001001001101011) && ({row_reg, col_reg}<20'b01100001010100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01100001010100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01100001010100011111) && ({row_reg, col_reg}<20'b01100001010101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01100001010101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01100001010101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01100001010101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01100001010101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01100001010101010000) && ({row_reg, col_reg}<20'b01100001011000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01100001011000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01100001011000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01100001011000111000) && ({row_reg, col_reg}<20'b01100001011000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01100001011000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01100001011000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01100001011000111100) && ({row_reg, col_reg}<20'b01100001011000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01100001011000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01100001011000111111) && ({row_reg, col_reg}<20'b01100001011001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01100001011001100110) && ({row_reg, col_reg}<20'b01100001011001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01100001011001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01100001011001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01100001011001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01100001011001101011) && ({row_reg, col_reg}<20'b01100001100100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01100001100100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01100001100100011111) && ({row_reg, col_reg}<20'b01100001100101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01100001100101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01100001100101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01100001100101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01100001100101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01100001100101010000) && ({row_reg, col_reg}<20'b01100001101000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01100001101000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01100001101000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01100001101000111000) && ({row_reg, col_reg}<20'b01100001101000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01100001101000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01100001101000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01100001101000111100) && ({row_reg, col_reg}<20'b01100001101000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01100001101000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01100001101000111111) && ({row_reg, col_reg}<20'b01100001101001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01100001101001100110) && ({row_reg, col_reg}<20'b01100001101001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01100001101001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01100001101001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01100001101001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01100001101001101011) && ({row_reg, col_reg}<20'b01100001110100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01100001110100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01100001110100011111) && ({row_reg, col_reg}<20'b01100001110101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01100001110101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01100001110101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01100001110101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01100001110101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01100001110101010000) && ({row_reg, col_reg}<20'b01100001111000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01100001111000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01100001111000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01100001111000111000) && ({row_reg, col_reg}<20'b01100001111000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01100001111000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01100001111000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01100001111000111100) && ({row_reg, col_reg}<20'b01100001111000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01100001111000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01100001111000111111) && ({row_reg, col_reg}<20'b01100001111001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01100001111001100110) && ({row_reg, col_reg}<20'b01100001111001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01100001111001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01100001111001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01100001111001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01100001111001101011) && ({row_reg, col_reg}<20'b01100010000100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01100010000100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01100010000100011111) && ({row_reg, col_reg}<20'b01100010000101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01100010000101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01100010000101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01100010000101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01100010000101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01100010000101010000) && ({row_reg, col_reg}<20'b01100010001000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01100010001000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01100010001000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01100010001000111000) && ({row_reg, col_reg}<20'b01100010001000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01100010001000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01100010001000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01100010001000111100) && ({row_reg, col_reg}<20'b01100010001000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01100010001000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01100010001000111111) && ({row_reg, col_reg}<20'b01100010001001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01100010001001100110) && ({row_reg, col_reg}<20'b01100010001001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01100010001001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01100010001001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01100010001001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01100010001001101011) && ({row_reg, col_reg}<20'b01100010010100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01100010010100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01100010010100011111) && ({row_reg, col_reg}<20'b01100010010101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01100010010101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01100010010101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01100010010101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01100010010101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01100010010101010000) && ({row_reg, col_reg}<20'b01100010011000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01100010011000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01100010011000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01100010011000111000) && ({row_reg, col_reg}<20'b01100010011000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01100010011000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01100010011000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01100010011000111100) && ({row_reg, col_reg}<20'b01100010011000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01100010011000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01100010011000111111) && ({row_reg, col_reg}<20'b01100010011001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01100010011001100110) && ({row_reg, col_reg}<20'b01100010011001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01100010011001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01100010011001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01100010011001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01100010011001101011) && ({row_reg, col_reg}<20'b01100010100100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01100010100100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01100010100100011111) && ({row_reg, col_reg}<20'b01100010100101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01100010100101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01100010100101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01100010100101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01100010100101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01100010100101010000) && ({row_reg, col_reg}<20'b01100010101000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01100010101000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01100010101000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01100010101000111000) && ({row_reg, col_reg}<20'b01100010101000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01100010101000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01100010101000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01100010101000111100) && ({row_reg, col_reg}<20'b01100010101000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01100010101000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01100010101000111111) && ({row_reg, col_reg}<20'b01100010101001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01100010101001100110) && ({row_reg, col_reg}<20'b01100010101001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01100010101001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01100010101001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01100010101001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01100010101001101011) && ({row_reg, col_reg}<20'b01100010110100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01100010110100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01100010110100011111) && ({row_reg, col_reg}<20'b01100010110101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01100010110101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01100010110101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01100010110101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01100010110101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01100010110101010000) && ({row_reg, col_reg}<20'b01100010111000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01100010111000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01100010111000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01100010111000111000) && ({row_reg, col_reg}<20'b01100010111000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01100010111000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01100010111000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01100010111000111100) && ({row_reg, col_reg}<20'b01100010111000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01100010111000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01100010111000111111) && ({row_reg, col_reg}<20'b01100010111001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01100010111001100110) && ({row_reg, col_reg}<20'b01100010111001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01100010111001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01100010111001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01100010111001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01100010111001101011) && ({row_reg, col_reg}<20'b01100011000100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01100011000100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01100011000100011111) && ({row_reg, col_reg}<20'b01100011000101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01100011000101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01100011000101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01100011000101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01100011000101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01100011000101010000) && ({row_reg, col_reg}<20'b01100011001000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01100011001000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01100011001000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01100011001000111000) && ({row_reg, col_reg}<20'b01100011001000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01100011001000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01100011001000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01100011001000111100) && ({row_reg, col_reg}<20'b01100011001000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01100011001000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01100011001000111111) && ({row_reg, col_reg}<20'b01100011001001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01100011001001100110) && ({row_reg, col_reg}<20'b01100011001001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01100011001001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01100011001001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01100011001001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01100011001001101011) && ({row_reg, col_reg}<20'b01100011010100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01100011010100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01100011010100011111) && ({row_reg, col_reg}<20'b01100011010101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01100011010101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01100011010101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01100011010101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01100011010101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01100011010101010000) && ({row_reg, col_reg}<20'b01100011011000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01100011011000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01100011011000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01100011011000111000) && ({row_reg, col_reg}<20'b01100011011000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01100011011000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01100011011000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01100011011000111100) && ({row_reg, col_reg}<20'b01100011011000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01100011011000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01100011011000111111) && ({row_reg, col_reg}<20'b01100011011001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01100011011001100110) && ({row_reg, col_reg}<20'b01100011011001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01100011011001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01100011011001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01100011011001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01100011011001101011) && ({row_reg, col_reg}<20'b01100011100100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01100011100100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01100011100100011111) && ({row_reg, col_reg}<20'b01100011100101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01100011100101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01100011100101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01100011100101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01100011100101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01100011100101010000) && ({row_reg, col_reg}<20'b01100011101000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01100011101000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01100011101000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01100011101000111000) && ({row_reg, col_reg}<20'b01100011101000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01100011101000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01100011101000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01100011101000111100) && ({row_reg, col_reg}<20'b01100011101000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01100011101000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01100011101000111111) && ({row_reg, col_reg}<20'b01100011101001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01100011101001100110) && ({row_reg, col_reg}<20'b01100011101001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01100011101001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01100011101001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01100011101001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01100011101001101011) && ({row_reg, col_reg}<20'b01100011110100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01100011110100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01100011110100011111) && ({row_reg, col_reg}<20'b01100011110101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01100011110101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01100011110101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01100011110101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01100011110101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01100011110101010000) && ({row_reg, col_reg}<20'b01100011111000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01100011111000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01100011111000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01100011111000111000) && ({row_reg, col_reg}<20'b01100011111000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01100011111000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01100011111000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01100011111000111100) && ({row_reg, col_reg}<20'b01100011111000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01100011111000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01100011111000111111) && ({row_reg, col_reg}<20'b01100011111001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01100011111001100110) && ({row_reg, col_reg}<20'b01100011111001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01100011111001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01100011111001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01100011111001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01100011111001101011) && ({row_reg, col_reg}<20'b01100100000100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01100100000100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01100100000100011111) && ({row_reg, col_reg}<20'b01100100000101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01100100000101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01100100000101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01100100000101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01100100000101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01100100000101010000) && ({row_reg, col_reg}<20'b01100100001000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01100100001000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01100100001000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01100100001000111000) && ({row_reg, col_reg}<20'b01100100001000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01100100001000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01100100001000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01100100001000111100) && ({row_reg, col_reg}<20'b01100100001000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01100100001000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01100100001000111111) && ({row_reg, col_reg}<20'b01100100001001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01100100001001100110) && ({row_reg, col_reg}<20'b01100100001001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01100100001001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01100100001001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01100100001001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01100100001001101011) && ({row_reg, col_reg}<20'b01100100010100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01100100010100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01100100010100011111) && ({row_reg, col_reg}<20'b01100100010101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01100100010101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01100100010101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01100100010101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01100100010101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01100100010101010000) && ({row_reg, col_reg}<20'b01100100011000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01100100011000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01100100011000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01100100011000111000) && ({row_reg, col_reg}<20'b01100100011000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01100100011000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01100100011000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01100100011000111100) && ({row_reg, col_reg}<20'b01100100011000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01100100011000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01100100011000111111) && ({row_reg, col_reg}<20'b01100100011001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01100100011001100110) && ({row_reg, col_reg}<20'b01100100011001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01100100011001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01100100011001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01100100011001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01100100011001101011) && ({row_reg, col_reg}<20'b01100100100100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01100100100100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01100100100100011111) && ({row_reg, col_reg}<20'b01100100100101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01100100100101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01100100100101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01100100100101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01100100100101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01100100100101010000) && ({row_reg, col_reg}<20'b01100100101000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01100100101000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01100100101000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01100100101000111000) && ({row_reg, col_reg}<20'b01100100101000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01100100101000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01100100101000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01100100101000111100) && ({row_reg, col_reg}<20'b01100100101000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01100100101000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01100100101000111111) && ({row_reg, col_reg}<20'b01100100101001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01100100101001100110) && ({row_reg, col_reg}<20'b01100100101001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01100100101001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01100100101001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01100100101001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01100100101001101011) && ({row_reg, col_reg}<20'b01100100110100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01100100110100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01100100110100011111) && ({row_reg, col_reg}<20'b01100100110101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01100100110101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01100100110101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01100100110101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01100100110101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01100100110101010000) && ({row_reg, col_reg}<20'b01100100111000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01100100111000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01100100111000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01100100111000111000) && ({row_reg, col_reg}<20'b01100100111000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01100100111000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01100100111000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01100100111000111100) && ({row_reg, col_reg}<20'b01100100111000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01100100111000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01100100111000111111) && ({row_reg, col_reg}<20'b01100100111001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01100100111001100110) && ({row_reg, col_reg}<20'b01100100111001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01100100111001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01100100111001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01100100111001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01100100111001101011) && ({row_reg, col_reg}<20'b01100101000100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01100101000100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01100101000100011111) && ({row_reg, col_reg}<20'b01100101000101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01100101000101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01100101000101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01100101000101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01100101000101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01100101000101010000) && ({row_reg, col_reg}<20'b01100101001000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01100101001000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01100101001000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01100101001000111000) && ({row_reg, col_reg}<20'b01100101001000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01100101001000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01100101001000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01100101001000111100) && ({row_reg, col_reg}<20'b01100101001000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01100101001000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01100101001000111111) && ({row_reg, col_reg}<20'b01100101001001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01100101001001100110) && ({row_reg, col_reg}<20'b01100101001001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01100101001001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01100101001001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01100101001001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01100101001001101011) && ({row_reg, col_reg}<20'b01100101010100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01100101010100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01100101010100011111) && ({row_reg, col_reg}<20'b01100101010101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01100101010101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01100101010101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01100101010101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01100101010101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01100101010101010000) && ({row_reg, col_reg}<20'b01100101011000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01100101011000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01100101011000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01100101011000111000) && ({row_reg, col_reg}<20'b01100101011000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01100101011000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01100101011000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01100101011000111100) && ({row_reg, col_reg}<20'b01100101011000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01100101011000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01100101011000111111) && ({row_reg, col_reg}<20'b01100101011001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01100101011001100110) && ({row_reg, col_reg}<20'b01100101011001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01100101011001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01100101011001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01100101011001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01100101011001101011) && ({row_reg, col_reg}<20'b01100101100100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01100101100100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01100101100100011111) && ({row_reg, col_reg}<20'b01100101100101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01100101100101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01100101100101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01100101100101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01100101100101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01100101100101010000) && ({row_reg, col_reg}<20'b01100101101000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01100101101000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01100101101000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01100101101000111000) && ({row_reg, col_reg}<20'b01100101101000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01100101101000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01100101101000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01100101101000111100) && ({row_reg, col_reg}<20'b01100101101000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01100101101000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01100101101000111111) && ({row_reg, col_reg}<20'b01100101101001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01100101101001100110) && ({row_reg, col_reg}<20'b01100101101001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01100101101001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01100101101001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01100101101001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01100101101001101011) && ({row_reg, col_reg}<20'b01100101110100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01100101110100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01100101110100011111) && ({row_reg, col_reg}<20'b01100101110101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01100101110101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01100101110101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01100101110101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01100101110101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01100101110101010000) && ({row_reg, col_reg}<20'b01100101111000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01100101111000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01100101111000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01100101111000111000) && ({row_reg, col_reg}<20'b01100101111000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01100101111000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01100101111000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01100101111000111100) && ({row_reg, col_reg}<20'b01100101111000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01100101111000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01100101111000111111) && ({row_reg, col_reg}<20'b01100101111001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01100101111001100110) && ({row_reg, col_reg}<20'b01100101111001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01100101111001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01100101111001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01100101111001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01100101111001101011) && ({row_reg, col_reg}<20'b01100110000100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01100110000100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01100110000100011111) && ({row_reg, col_reg}<20'b01100110000101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01100110000101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01100110000101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01100110000101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01100110000101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01100110000101010000) && ({row_reg, col_reg}<20'b01100110001000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01100110001000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01100110001000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01100110001000111000) && ({row_reg, col_reg}<20'b01100110001000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01100110001000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01100110001000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01100110001000111100) && ({row_reg, col_reg}<20'b01100110001000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01100110001000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01100110001000111111) && ({row_reg, col_reg}<20'b01100110001001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01100110001001100110) && ({row_reg, col_reg}<20'b01100110001001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01100110001001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01100110001001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01100110001001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01100110001001101011) && ({row_reg, col_reg}<20'b01100110010100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01100110010100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01100110010100011111) && ({row_reg, col_reg}<20'b01100110010101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01100110010101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01100110010101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01100110010101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01100110010101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01100110010101010000) && ({row_reg, col_reg}<20'b01100110011000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01100110011000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01100110011000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01100110011000111000) && ({row_reg, col_reg}<20'b01100110011000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01100110011000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01100110011000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01100110011000111100) && ({row_reg, col_reg}<20'b01100110011000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01100110011000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01100110011000111111) && ({row_reg, col_reg}<20'b01100110011001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01100110011001100110) && ({row_reg, col_reg}<20'b01100110011001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01100110011001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01100110011001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01100110011001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01100110011001101011) && ({row_reg, col_reg}<20'b01100110100100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01100110100100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01100110100100011111) && ({row_reg, col_reg}<20'b01100110100101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01100110100101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01100110100101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01100110100101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01100110100101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01100110100101010000) && ({row_reg, col_reg}<20'b01100110101000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01100110101000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01100110101000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01100110101000111000) && ({row_reg, col_reg}<20'b01100110101000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01100110101000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01100110101000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01100110101000111100) && ({row_reg, col_reg}<20'b01100110101000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01100110101000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01100110101000111111) && ({row_reg, col_reg}<20'b01100110101001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01100110101001100110) && ({row_reg, col_reg}<20'b01100110101001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01100110101001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01100110101001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01100110101001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01100110101001101011) && ({row_reg, col_reg}<20'b01100110110100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01100110110100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01100110110100011111) && ({row_reg, col_reg}<20'b01100110110101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01100110110101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01100110110101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01100110110101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01100110110101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01100110110101010000) && ({row_reg, col_reg}<20'b01100110111000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01100110111000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01100110111000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01100110111000111000) && ({row_reg, col_reg}<20'b01100110111000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01100110111000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01100110111000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01100110111000111100) && ({row_reg, col_reg}<20'b01100110111000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01100110111000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01100110111000111111) && ({row_reg, col_reg}<20'b01100110111001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01100110111001100110) && ({row_reg, col_reg}<20'b01100110111001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01100110111001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01100110111001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01100110111001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01100110111001101011) && ({row_reg, col_reg}<20'b01100111000100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01100111000100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01100111000100011111) && ({row_reg, col_reg}<20'b01100111000101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01100111000101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01100111000101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01100111000101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01100111000101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01100111000101010000) && ({row_reg, col_reg}<20'b01100111001000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01100111001000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01100111001000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01100111001000111000) && ({row_reg, col_reg}<20'b01100111001000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01100111001000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01100111001000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01100111001000111100) && ({row_reg, col_reg}<20'b01100111001000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01100111001000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01100111001000111111) && ({row_reg, col_reg}<20'b01100111001001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01100111001001100110) && ({row_reg, col_reg}<20'b01100111001001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01100111001001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01100111001001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01100111001001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01100111001001101011) && ({row_reg, col_reg}<20'b01100111010100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01100111010100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01100111010100011111) && ({row_reg, col_reg}<20'b01100111010101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01100111010101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01100111010101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01100111010101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01100111010101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01100111010101010000) && ({row_reg, col_reg}<20'b01100111011000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01100111011000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01100111011000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01100111011000111000) && ({row_reg, col_reg}<20'b01100111011000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01100111011000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01100111011000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01100111011000111100) && ({row_reg, col_reg}<20'b01100111011000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01100111011000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01100111011000111111) && ({row_reg, col_reg}<20'b01100111011001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01100111011001100110) && ({row_reg, col_reg}<20'b01100111011001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01100111011001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01100111011001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01100111011001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01100111011001101011) && ({row_reg, col_reg}<20'b01100111100100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01100111100100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01100111100100011111) && ({row_reg, col_reg}<20'b01100111100101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01100111100101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01100111100101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01100111100101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01100111100101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01100111100101010000) && ({row_reg, col_reg}<20'b01100111101000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01100111101000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01100111101000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01100111101000111000) && ({row_reg, col_reg}<20'b01100111101000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01100111101000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01100111101000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01100111101000111100) && ({row_reg, col_reg}<20'b01100111101000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01100111101000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01100111101000111111) && ({row_reg, col_reg}<20'b01100111101001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01100111101001100110) && ({row_reg, col_reg}<20'b01100111101001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01100111101001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01100111101001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01100111101001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01100111101001101011) && ({row_reg, col_reg}<20'b01100111110100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01100111110100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01100111110100011111) && ({row_reg, col_reg}<20'b01100111110101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01100111110101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01100111110101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01100111110101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01100111110101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01100111110101010000) && ({row_reg, col_reg}<20'b01100111111000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01100111111000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01100111111000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01100111111000111000) && ({row_reg, col_reg}<20'b01100111111000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01100111111000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01100111111000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01100111111000111100) && ({row_reg, col_reg}<20'b01100111111000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01100111111000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01100111111000111111) && ({row_reg, col_reg}<20'b01100111111001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01100111111001100110) && ({row_reg, col_reg}<20'b01100111111001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01100111111001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01100111111001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01100111111001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01100111111001101011) && ({row_reg, col_reg}<20'b01101000000100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01101000000100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01101000000100011111) && ({row_reg, col_reg}<20'b01101000000101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01101000000101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01101000000101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01101000000101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01101000000101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01101000000101010000) && ({row_reg, col_reg}<20'b01101000001000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01101000001000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01101000001000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01101000001000111000) && ({row_reg, col_reg}<20'b01101000001000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01101000001000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01101000001000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01101000001000111100) && ({row_reg, col_reg}<20'b01101000001000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01101000001000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01101000001000111111) && ({row_reg, col_reg}<20'b01101000001001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01101000001001100110) && ({row_reg, col_reg}<20'b01101000001001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01101000001001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01101000001001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01101000001001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01101000001001101011) && ({row_reg, col_reg}<20'b01101000010100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01101000010100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01101000010100011111) && ({row_reg, col_reg}<20'b01101000010101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01101000010101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01101000010101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01101000010101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01101000010101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01101000010101010000) && ({row_reg, col_reg}<20'b01101000011000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01101000011000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01101000011000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01101000011000111000) && ({row_reg, col_reg}<20'b01101000011000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01101000011000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01101000011000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01101000011000111100) && ({row_reg, col_reg}<20'b01101000011000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01101000011000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01101000011000111111) && ({row_reg, col_reg}<20'b01101000011001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01101000011001100110) && ({row_reg, col_reg}<20'b01101000011001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01101000011001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01101000011001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01101000011001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01101000011001101011) && ({row_reg, col_reg}<20'b01101000100100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01101000100100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01101000100100011111) && ({row_reg, col_reg}<20'b01101000100101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01101000100101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01101000100101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01101000100101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01101000100101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01101000100101010000) && ({row_reg, col_reg}<20'b01101000101000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01101000101000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01101000101000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01101000101000111000) && ({row_reg, col_reg}<20'b01101000101000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01101000101000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01101000101000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01101000101000111100) && ({row_reg, col_reg}<20'b01101000101000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01101000101000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01101000101000111111) && ({row_reg, col_reg}<20'b01101000101001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01101000101001100110) && ({row_reg, col_reg}<20'b01101000101001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01101000101001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01101000101001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01101000101001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01101000101001101011) && ({row_reg, col_reg}<20'b01101000110100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01101000110100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01101000110100011111) && ({row_reg, col_reg}<20'b01101000110101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01101000110101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01101000110101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01101000110101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01101000110101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01101000110101010000) && ({row_reg, col_reg}<20'b01101000111000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01101000111000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01101000111000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01101000111000111000) && ({row_reg, col_reg}<20'b01101000111000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01101000111000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01101000111000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01101000111000111100) && ({row_reg, col_reg}<20'b01101000111000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01101000111000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01101000111000111111) && ({row_reg, col_reg}<20'b01101000111001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01101000111001100110) && ({row_reg, col_reg}<20'b01101000111001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01101000111001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01101000111001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01101000111001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01101000111001101011) && ({row_reg, col_reg}<20'b01101001000100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01101001000100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01101001000100011111) && ({row_reg, col_reg}<20'b01101001000101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01101001000101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01101001000101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01101001000101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01101001000101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01101001000101010000) && ({row_reg, col_reg}<20'b01101001001000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01101001001000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01101001001000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01101001001000111000) && ({row_reg, col_reg}<20'b01101001001000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01101001001000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01101001001000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01101001001000111100) && ({row_reg, col_reg}<20'b01101001001000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01101001001000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01101001001000111111) && ({row_reg, col_reg}<20'b01101001001001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01101001001001100110) && ({row_reg, col_reg}<20'b01101001001001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01101001001001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01101001001001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01101001001001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01101001001001101011) && ({row_reg, col_reg}<20'b01101001010100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01101001010100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01101001010100011111) && ({row_reg, col_reg}<20'b01101001010101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01101001010101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01101001010101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01101001010101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01101001010101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01101001010101010000) && ({row_reg, col_reg}<20'b01101001011000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01101001011000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01101001011000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01101001011000111000) && ({row_reg, col_reg}<20'b01101001011000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01101001011000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01101001011000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01101001011000111100) && ({row_reg, col_reg}<20'b01101001011000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01101001011000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01101001011000111111) && ({row_reg, col_reg}<20'b01101001011001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01101001011001100110) && ({row_reg, col_reg}<20'b01101001011001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01101001011001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01101001011001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01101001011001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01101001011001101011) && ({row_reg, col_reg}<20'b01101001100100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01101001100100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01101001100100011111) && ({row_reg, col_reg}<20'b01101001100101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01101001100101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01101001100101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01101001100101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01101001100101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01101001100101010000) && ({row_reg, col_reg}<20'b01101001101000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01101001101000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01101001101000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01101001101000111000) && ({row_reg, col_reg}<20'b01101001101000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01101001101000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01101001101000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01101001101000111100) && ({row_reg, col_reg}<20'b01101001101000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01101001101000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01101001101000111111) && ({row_reg, col_reg}<20'b01101001101001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01101001101001100110) && ({row_reg, col_reg}<20'b01101001101001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01101001101001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01101001101001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01101001101001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01101001101001101011) && ({row_reg, col_reg}<20'b01101001110100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01101001110100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01101001110100011111) && ({row_reg, col_reg}<20'b01101001110101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01101001110101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01101001110101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01101001110101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01101001110101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01101001110101010000) && ({row_reg, col_reg}<20'b01101001111000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01101001111000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01101001111000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01101001111000111000) && ({row_reg, col_reg}<20'b01101001111000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01101001111000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01101001111000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01101001111000111100) && ({row_reg, col_reg}<20'b01101001111000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01101001111000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01101001111000111111) && ({row_reg, col_reg}<20'b01101001111001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01101001111001100110) && ({row_reg, col_reg}<20'b01101001111001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01101001111001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01101001111001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01101001111001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01101001111001101011) && ({row_reg, col_reg}<20'b01101010000100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01101010000100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01101010000100011111) && ({row_reg, col_reg}<20'b01101010000101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01101010000101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01101010000101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01101010000101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01101010000101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01101010000101010000) && ({row_reg, col_reg}<20'b01101010001000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01101010001000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01101010001000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01101010001000111000) && ({row_reg, col_reg}<20'b01101010001000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01101010001000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01101010001000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01101010001000111100) && ({row_reg, col_reg}<20'b01101010001000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01101010001000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01101010001000111111) && ({row_reg, col_reg}<20'b01101010001001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01101010001001100110) && ({row_reg, col_reg}<20'b01101010001001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01101010001001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01101010001001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01101010001001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01101010001001101011) && ({row_reg, col_reg}<20'b01101010010100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01101010010100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01101010010100011111) && ({row_reg, col_reg}<20'b01101010010101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01101010010101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01101010010101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01101010010101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01101010010101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01101010010101010000) && ({row_reg, col_reg}<20'b01101010011000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01101010011000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01101010011000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01101010011000111000) && ({row_reg, col_reg}<20'b01101010011000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01101010011000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01101010011000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01101010011000111100) && ({row_reg, col_reg}<20'b01101010011000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01101010011000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01101010011000111111) && ({row_reg, col_reg}<20'b01101010011001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01101010011001100110) && ({row_reg, col_reg}<20'b01101010011001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01101010011001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01101010011001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01101010011001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01101010011001101011) && ({row_reg, col_reg}<20'b01101010100100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01101010100100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01101010100100011111) && ({row_reg, col_reg}<20'b01101010100101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01101010100101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01101010100101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01101010100101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01101010100101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01101010100101010000) && ({row_reg, col_reg}<20'b01101010101000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01101010101000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01101010101000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01101010101000111000) && ({row_reg, col_reg}<20'b01101010101000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01101010101000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01101010101000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01101010101000111100) && ({row_reg, col_reg}<20'b01101010101000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01101010101000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01101010101000111111) && ({row_reg, col_reg}<20'b01101010101001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01101010101001100110) && ({row_reg, col_reg}<20'b01101010101001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01101010101001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01101010101001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01101010101001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01101010101001101011) && ({row_reg, col_reg}<20'b01101010110100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01101010110100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01101010110100011111) && ({row_reg, col_reg}<20'b01101010110101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01101010110101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01101010110101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01101010110101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01101010110101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01101010110101010000) && ({row_reg, col_reg}<20'b01101010111000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01101010111000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01101010111000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01101010111000111000) && ({row_reg, col_reg}<20'b01101010111000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01101010111000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01101010111000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01101010111000111100) && ({row_reg, col_reg}<20'b01101010111000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01101010111000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01101010111000111111) && ({row_reg, col_reg}<20'b01101010111001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01101010111001100110) && ({row_reg, col_reg}<20'b01101010111001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01101010111001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01101010111001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01101010111001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01101010111001101011) && ({row_reg, col_reg}<20'b01101011000100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01101011000100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01101011000100011111) && ({row_reg, col_reg}<20'b01101011000101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01101011000101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01101011000101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01101011000101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01101011000101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01101011000101010000) && ({row_reg, col_reg}<20'b01101011001000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01101011001000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01101011001000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01101011001000111000) && ({row_reg, col_reg}<20'b01101011001000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01101011001000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01101011001000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01101011001000111100) && ({row_reg, col_reg}<20'b01101011001000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01101011001000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01101011001000111111) && ({row_reg, col_reg}<20'b01101011001001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01101011001001100110) && ({row_reg, col_reg}<20'b01101011001001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01101011001001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01101011001001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01101011001001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01101011001001101011) && ({row_reg, col_reg}<20'b01101011010100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01101011010100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01101011010100011111) && ({row_reg, col_reg}<20'b01101011010101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01101011010101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01101011010101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01101011010101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01101011010101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01101011010101010000) && ({row_reg, col_reg}<20'b01101011011000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01101011011000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01101011011000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01101011011000111000) && ({row_reg, col_reg}<20'b01101011011000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01101011011000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01101011011000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01101011011000111100) && ({row_reg, col_reg}<20'b01101011011000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01101011011000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01101011011000111111) && ({row_reg, col_reg}<20'b01101011011001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01101011011001100110) && ({row_reg, col_reg}<20'b01101011011001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01101011011001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01101011011001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01101011011001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01101011011001101011) && ({row_reg, col_reg}<20'b01101011100100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01101011100100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01101011100100011111) && ({row_reg, col_reg}<20'b01101011100101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01101011100101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01101011100101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01101011100101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01101011100101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01101011100101010000) && ({row_reg, col_reg}<20'b01101011101000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01101011101000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01101011101000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01101011101000111000) && ({row_reg, col_reg}<20'b01101011101000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01101011101000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01101011101000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01101011101000111100) && ({row_reg, col_reg}<20'b01101011101000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01101011101000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01101011101000111111) && ({row_reg, col_reg}<20'b01101011101001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01101011101001100110) && ({row_reg, col_reg}<20'b01101011101001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01101011101001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01101011101001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01101011101001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01101011101001101011) && ({row_reg, col_reg}<20'b01101011110100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01101011110100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01101011110100011111) && ({row_reg, col_reg}<20'b01101011110101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01101011110101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01101011110101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01101011110101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01101011110101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01101011110101010000) && ({row_reg, col_reg}<20'b01101011111000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01101011111000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01101011111000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01101011111000111000) && ({row_reg, col_reg}<20'b01101011111000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01101011111000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01101011111000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01101011111000111100) && ({row_reg, col_reg}<20'b01101011111000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01101011111000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01101011111000111111) && ({row_reg, col_reg}<20'b01101011111001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01101011111001100110) && ({row_reg, col_reg}<20'b01101011111001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01101011111001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01101011111001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01101011111001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01101011111001101011) && ({row_reg, col_reg}<20'b01101100000100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01101100000100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01101100000100011111) && ({row_reg, col_reg}<20'b01101100000101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01101100000101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01101100000101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01101100000101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01101100000101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01101100000101010000) && ({row_reg, col_reg}<20'b01101100001000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01101100001000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01101100001000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01101100001000111000) && ({row_reg, col_reg}<20'b01101100001000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01101100001000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01101100001000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01101100001000111100) && ({row_reg, col_reg}<20'b01101100001000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01101100001000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01101100001000111111) && ({row_reg, col_reg}<20'b01101100001001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01101100001001100110) && ({row_reg, col_reg}<20'b01101100001001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01101100001001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01101100001001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01101100001001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01101100001001101011) && ({row_reg, col_reg}<20'b01101100010100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01101100010100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01101100010100011111) && ({row_reg, col_reg}<20'b01101100010101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01101100010101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01101100010101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01101100010101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01101100010101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01101100010101010000) && ({row_reg, col_reg}<20'b01101100011000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01101100011000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01101100011000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01101100011000111000) && ({row_reg, col_reg}<20'b01101100011000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01101100011000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01101100011000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01101100011000111100) && ({row_reg, col_reg}<20'b01101100011000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01101100011000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01101100011000111111) && ({row_reg, col_reg}<20'b01101100011001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01101100011001100110) && ({row_reg, col_reg}<20'b01101100011001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01101100011001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01101100011001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01101100011001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01101100011001101011) && ({row_reg, col_reg}<20'b01101100100100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01101100100100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01101100100100011111) && ({row_reg, col_reg}<20'b01101100100101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01101100100101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01101100100101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01101100100101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01101100100101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01101100100101010000) && ({row_reg, col_reg}<20'b01101100101000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01101100101000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01101100101000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01101100101000111000) && ({row_reg, col_reg}<20'b01101100101000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01101100101000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01101100101000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01101100101000111100) && ({row_reg, col_reg}<20'b01101100101000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01101100101000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01101100101000111111) && ({row_reg, col_reg}<20'b01101100101001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01101100101001100110) && ({row_reg, col_reg}<20'b01101100101001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01101100101001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01101100101001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01101100101001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01101100101001101011) && ({row_reg, col_reg}<20'b01101100110100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01101100110100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01101100110100011111) && ({row_reg, col_reg}<20'b01101100110101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01101100110101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01101100110101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01101100110101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01101100110101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01101100110101010000) && ({row_reg, col_reg}<20'b01101100111000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01101100111000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01101100111000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01101100111000111000) && ({row_reg, col_reg}<20'b01101100111000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01101100111000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01101100111000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01101100111000111100) && ({row_reg, col_reg}<20'b01101100111000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01101100111000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01101100111000111111) && ({row_reg, col_reg}<20'b01101100111001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01101100111001100110) && ({row_reg, col_reg}<20'b01101100111001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01101100111001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01101100111001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01101100111001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01101100111001101011) && ({row_reg, col_reg}<20'b01101101000100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01101101000100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01101101000100011111) && ({row_reg, col_reg}<20'b01101101000101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01101101000101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01101101000101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01101101000101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01101101000101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01101101000101010000) && ({row_reg, col_reg}<20'b01101101001000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01101101001000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01101101001000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01101101001000111000) && ({row_reg, col_reg}<20'b01101101001000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01101101001000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01101101001000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01101101001000111100) && ({row_reg, col_reg}<20'b01101101001000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01101101001000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01101101001000111111) && ({row_reg, col_reg}<20'b01101101001001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01101101001001100110) && ({row_reg, col_reg}<20'b01101101001001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01101101001001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01101101001001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01101101001001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01101101001001101011) && ({row_reg, col_reg}<20'b01101101010100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01101101010100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01101101010100011111) && ({row_reg, col_reg}<20'b01101101010101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01101101010101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01101101010101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01101101010101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01101101010101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01101101010101010000) && ({row_reg, col_reg}<20'b01101101011000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01101101011000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01101101011000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01101101011000111000) && ({row_reg, col_reg}<20'b01101101011000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01101101011000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01101101011000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01101101011000111100) && ({row_reg, col_reg}<20'b01101101011000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01101101011000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01101101011000111111) && ({row_reg, col_reg}<20'b01101101011001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01101101011001100110) && ({row_reg, col_reg}<20'b01101101011001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01101101011001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01101101011001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01101101011001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01101101011001101011) && ({row_reg, col_reg}<20'b01101101100100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01101101100100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01101101100100011111) && ({row_reg, col_reg}<20'b01101101100101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01101101100101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01101101100101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01101101100101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01101101100101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01101101100101010000) && ({row_reg, col_reg}<20'b01101101101000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01101101101000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01101101101000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01101101101000111000) && ({row_reg, col_reg}<20'b01101101101000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01101101101000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01101101101000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01101101101000111100) && ({row_reg, col_reg}<20'b01101101101000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01101101101000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01101101101000111111) && ({row_reg, col_reg}<20'b01101101101001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01101101101001100110) && ({row_reg, col_reg}<20'b01101101101001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01101101101001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01101101101001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01101101101001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01101101101001101011) && ({row_reg, col_reg}<20'b01101101110100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01101101110100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01101101110100011111) && ({row_reg, col_reg}<20'b01101101110101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01101101110101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01101101110101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01101101110101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01101101110101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01101101110101010000) && ({row_reg, col_reg}<20'b01101101111000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01101101111000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01101101111000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01101101111000111000) && ({row_reg, col_reg}<20'b01101101111000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01101101111000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01101101111000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01101101111000111100) && ({row_reg, col_reg}<20'b01101101111000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01101101111000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01101101111000111111) && ({row_reg, col_reg}<20'b01101101111001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01101101111001100110) && ({row_reg, col_reg}<20'b01101101111001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01101101111001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01101101111001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01101101111001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01101101111001101011) && ({row_reg, col_reg}<20'b01101110000100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01101110000100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01101110000100011111) && ({row_reg, col_reg}<20'b01101110000101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01101110000101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01101110000101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01101110000101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01101110000101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01101110000101010000) && ({row_reg, col_reg}<20'b01101110001000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01101110001000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01101110001000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01101110001000111000) && ({row_reg, col_reg}<20'b01101110001000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01101110001000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01101110001000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01101110001000111100) && ({row_reg, col_reg}<20'b01101110001000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01101110001000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01101110001000111111) && ({row_reg, col_reg}<20'b01101110001001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01101110001001100110) && ({row_reg, col_reg}<20'b01101110001001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01101110001001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01101110001001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01101110001001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01101110001001101011) && ({row_reg, col_reg}<20'b01101110010100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01101110010100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01101110010100011111) && ({row_reg, col_reg}<20'b01101110010101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01101110010101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01101110010101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01101110010101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01101110010101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01101110010101010000) && ({row_reg, col_reg}<20'b01101110011000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01101110011000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01101110011000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01101110011000111000) && ({row_reg, col_reg}<20'b01101110011000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01101110011000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01101110011000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01101110011000111100) && ({row_reg, col_reg}<20'b01101110011000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01101110011000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01101110011000111111) && ({row_reg, col_reg}<20'b01101110011001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01101110011001100110) && ({row_reg, col_reg}<20'b01101110011001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01101110011001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01101110011001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01101110011001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01101110011001101011) && ({row_reg, col_reg}<20'b01101110100100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01101110100100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01101110100100011111) && ({row_reg, col_reg}<20'b01101110100101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01101110100101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01101110100101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01101110100101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01101110100101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01101110100101010000) && ({row_reg, col_reg}<20'b01101110101000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01101110101000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01101110101000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01101110101000111000) && ({row_reg, col_reg}<20'b01101110101000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01101110101000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01101110101000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01101110101000111100) && ({row_reg, col_reg}<20'b01101110101000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01101110101000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01101110101000111111) && ({row_reg, col_reg}<20'b01101110101001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01101110101001100110) && ({row_reg, col_reg}<20'b01101110101001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01101110101001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01101110101001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01101110101001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01101110101001101011) && ({row_reg, col_reg}<20'b01101110110100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01101110110100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01101110110100011111) && ({row_reg, col_reg}<20'b01101110110101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01101110110101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01101110110101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01101110110101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01101110110101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01101110110101010000) && ({row_reg, col_reg}<20'b01101110111000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01101110111000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01101110111000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01101110111000111000) && ({row_reg, col_reg}<20'b01101110111000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01101110111000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01101110111000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01101110111000111100) && ({row_reg, col_reg}<20'b01101110111000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01101110111000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01101110111000111111) && ({row_reg, col_reg}<20'b01101110111001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01101110111001100110) && ({row_reg, col_reg}<20'b01101110111001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01101110111001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01101110111001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01101110111001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01101110111001101011) && ({row_reg, col_reg}<20'b01101111000100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01101111000100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01101111000100011111) && ({row_reg, col_reg}<20'b01101111000101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01101111000101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01101111000101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01101111000101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01101111000101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01101111000101010000) && ({row_reg, col_reg}<20'b01101111001000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01101111001000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01101111001000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01101111001000111000) && ({row_reg, col_reg}<20'b01101111001000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01101111001000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01101111001000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01101111001000111100) && ({row_reg, col_reg}<20'b01101111001000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01101111001000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01101111001000111111) && ({row_reg, col_reg}<20'b01101111001001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01101111001001100110) && ({row_reg, col_reg}<20'b01101111001001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01101111001001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01101111001001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01101111001001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01101111001001101011) && ({row_reg, col_reg}<20'b01101111010100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01101111010100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01101111010100011111) && ({row_reg, col_reg}<20'b01101111010101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01101111010101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01101111010101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01101111010101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01101111010101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01101111010101010000) && ({row_reg, col_reg}<20'b01101111011000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01101111011000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01101111011000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01101111011000111000) && ({row_reg, col_reg}<20'b01101111011000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01101111011000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01101111011000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01101111011000111100) && ({row_reg, col_reg}<20'b01101111011000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01101111011000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01101111011000111111) && ({row_reg, col_reg}<20'b01101111011001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01101111011001100110) && ({row_reg, col_reg}<20'b01101111011001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01101111011001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01101111011001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01101111011001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01101111011001101011) && ({row_reg, col_reg}<20'b01101111100100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01101111100100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01101111100100011111) && ({row_reg, col_reg}<20'b01101111100101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01101111100101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01101111100101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01101111100101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01101111100101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01101111100101010000) && ({row_reg, col_reg}<20'b01101111101000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01101111101000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01101111101000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01101111101000111000) && ({row_reg, col_reg}<20'b01101111101000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01101111101000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01101111101000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01101111101000111100) && ({row_reg, col_reg}<20'b01101111101000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01101111101000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01101111101000111111) && ({row_reg, col_reg}<20'b01101111101001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01101111101001100110) && ({row_reg, col_reg}<20'b01101111101001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01101111101001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01101111101001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01101111101001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01101111101001101011) && ({row_reg, col_reg}<20'b01101111110100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01101111110100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01101111110100011111) && ({row_reg, col_reg}<20'b01101111110101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01101111110101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01101111110101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01101111110101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01101111110101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01101111110101010000) && ({row_reg, col_reg}<20'b01101111111000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01101111111000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01101111111000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01101111111000111000) && ({row_reg, col_reg}<20'b01101111111000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01101111111000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01101111111000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01101111111000111100) && ({row_reg, col_reg}<20'b01101111111000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01101111111000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01101111111000111111) && ({row_reg, col_reg}<20'b01101111111001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01101111111001100110) && ({row_reg, col_reg}<20'b01101111111001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01101111111001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01101111111001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01101111111001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01101111111001101011) && ({row_reg, col_reg}<20'b01110000000100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01110000000100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01110000000100011111) && ({row_reg, col_reg}<20'b01110000000101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01110000000101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01110000000101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01110000000101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01110000000101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01110000000101010000) && ({row_reg, col_reg}<20'b01110000001000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01110000001000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01110000001000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01110000001000111000) && ({row_reg, col_reg}<20'b01110000001000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01110000001000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01110000001000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01110000001000111100) && ({row_reg, col_reg}<20'b01110000001000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01110000001000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01110000001000111111) && ({row_reg, col_reg}<20'b01110000001001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01110000001001100110) && ({row_reg, col_reg}<20'b01110000001001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01110000001001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01110000001001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01110000001001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01110000001001101011) && ({row_reg, col_reg}<20'b01110000010100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01110000010100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01110000010100011111) && ({row_reg, col_reg}<20'b01110000010101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01110000010101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01110000010101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01110000010101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01110000010101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01110000010101010000) && ({row_reg, col_reg}<20'b01110000011000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01110000011000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01110000011000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01110000011000111000) && ({row_reg, col_reg}<20'b01110000011000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01110000011000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01110000011000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01110000011000111100) && ({row_reg, col_reg}<20'b01110000011000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01110000011000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01110000011000111111) && ({row_reg, col_reg}<20'b01110000011001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01110000011001100110) && ({row_reg, col_reg}<20'b01110000011001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01110000011001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01110000011001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01110000011001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01110000011001101011) && ({row_reg, col_reg}<20'b01110000100100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01110000100100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01110000100100011111) && ({row_reg, col_reg}<20'b01110000100101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01110000100101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01110000100101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01110000100101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01110000100101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01110000100101010000) && ({row_reg, col_reg}<20'b01110000101000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01110000101000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01110000101000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01110000101000111000) && ({row_reg, col_reg}<20'b01110000101000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01110000101000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01110000101000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01110000101000111100) && ({row_reg, col_reg}<20'b01110000101000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01110000101000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01110000101000111111) && ({row_reg, col_reg}<20'b01110000101001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01110000101001100110) && ({row_reg, col_reg}<20'b01110000101001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01110000101001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01110000101001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01110000101001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01110000101001101011) && ({row_reg, col_reg}<20'b01110000110100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01110000110100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01110000110100011111) && ({row_reg, col_reg}<20'b01110000110101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01110000110101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01110000110101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01110000110101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01110000110101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01110000110101010000) && ({row_reg, col_reg}<20'b01110000111000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01110000111000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01110000111000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01110000111000111000) && ({row_reg, col_reg}<20'b01110000111000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01110000111000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01110000111000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01110000111000111100) && ({row_reg, col_reg}<20'b01110000111000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01110000111000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01110000111000111111) && ({row_reg, col_reg}<20'b01110000111001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01110000111001100110) && ({row_reg, col_reg}<20'b01110000111001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01110000111001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01110000111001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01110000111001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01110000111001101011) && ({row_reg, col_reg}<20'b01110001000100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01110001000100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01110001000100011111) && ({row_reg, col_reg}<20'b01110001000101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01110001000101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01110001000101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01110001000101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01110001000101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01110001000101010000) && ({row_reg, col_reg}<20'b01110001001000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01110001001000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01110001001000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01110001001000111000) && ({row_reg, col_reg}<20'b01110001001000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01110001001000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01110001001000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01110001001000111100) && ({row_reg, col_reg}<20'b01110001001000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01110001001000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01110001001000111111) && ({row_reg, col_reg}<20'b01110001001001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01110001001001100110) && ({row_reg, col_reg}<20'b01110001001001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01110001001001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01110001001001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01110001001001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01110001001001101011) && ({row_reg, col_reg}<20'b01110001010100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01110001010100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01110001010100011111) && ({row_reg, col_reg}<20'b01110001010101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01110001010101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01110001010101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01110001010101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01110001010101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01110001010101010000) && ({row_reg, col_reg}<20'b01110001011000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01110001011000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01110001011000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01110001011000111000) && ({row_reg, col_reg}<20'b01110001011000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01110001011000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01110001011000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01110001011000111100) && ({row_reg, col_reg}<20'b01110001011000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01110001011000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01110001011000111111) && ({row_reg, col_reg}<20'b01110001011001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01110001011001100110) && ({row_reg, col_reg}<20'b01110001011001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01110001011001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01110001011001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01110001011001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01110001011001101011) && ({row_reg, col_reg}<20'b01110001100100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01110001100100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01110001100100011111) && ({row_reg, col_reg}<20'b01110001100101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01110001100101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01110001100101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01110001100101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01110001100101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01110001100101010000) && ({row_reg, col_reg}<20'b01110001101000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01110001101000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01110001101000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01110001101000111000) && ({row_reg, col_reg}<20'b01110001101000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01110001101000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01110001101000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01110001101000111100) && ({row_reg, col_reg}<20'b01110001101000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01110001101000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01110001101000111111) && ({row_reg, col_reg}<20'b01110001101001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01110001101001100110) && ({row_reg, col_reg}<20'b01110001101001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01110001101001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01110001101001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01110001101001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01110001101001101011) && ({row_reg, col_reg}<20'b01110001110100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01110001110100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01110001110100011111) && ({row_reg, col_reg}<20'b01110001110101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01110001110101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01110001110101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01110001110101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01110001110101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01110001110101010000) && ({row_reg, col_reg}<20'b01110001111000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01110001111000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01110001111000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01110001111000111000) && ({row_reg, col_reg}<20'b01110001111000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01110001111000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01110001111000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01110001111000111100) && ({row_reg, col_reg}<20'b01110001111000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01110001111000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01110001111000111111) && ({row_reg, col_reg}<20'b01110001111001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01110001111001100110) && ({row_reg, col_reg}<20'b01110001111001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01110001111001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01110001111001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01110001111001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01110001111001101011) && ({row_reg, col_reg}<20'b01110010000100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01110010000100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01110010000100011111) && ({row_reg, col_reg}<20'b01110010000101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01110010000101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01110010000101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01110010000101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01110010000101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01110010000101010000) && ({row_reg, col_reg}<20'b01110010001000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01110010001000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01110010001000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01110010001000111000) && ({row_reg, col_reg}<20'b01110010001000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01110010001000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01110010001000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01110010001000111100) && ({row_reg, col_reg}<20'b01110010001000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01110010001000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01110010001000111111) && ({row_reg, col_reg}<20'b01110010001001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01110010001001100110) && ({row_reg, col_reg}<20'b01110010001001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01110010001001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01110010001001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01110010001001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01110010001001101011) && ({row_reg, col_reg}<20'b01110010010100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01110010010100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01110010010100011111) && ({row_reg, col_reg}<20'b01110010010101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01110010010101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01110010010101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01110010010101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01110010010101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01110010010101010000) && ({row_reg, col_reg}<20'b01110010011000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01110010011000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01110010011000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01110010011000111000) && ({row_reg, col_reg}<20'b01110010011000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01110010011000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01110010011000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01110010011000111100) && ({row_reg, col_reg}<20'b01110010011000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01110010011000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01110010011000111111) && ({row_reg, col_reg}<20'b01110010011001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01110010011001100110) && ({row_reg, col_reg}<20'b01110010011001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01110010011001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01110010011001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01110010011001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01110010011001101011) && ({row_reg, col_reg}<20'b01110010100100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01110010100100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01110010100100011111) && ({row_reg, col_reg}<20'b01110010100101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01110010100101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01110010100101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01110010100101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01110010100101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01110010100101010000) && ({row_reg, col_reg}<20'b01110010101000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01110010101000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01110010101000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01110010101000111000) && ({row_reg, col_reg}<20'b01110010101000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01110010101000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01110010101000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01110010101000111100) && ({row_reg, col_reg}<20'b01110010101000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01110010101000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01110010101000111111) && ({row_reg, col_reg}<20'b01110010101001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01110010101001100110) && ({row_reg, col_reg}<20'b01110010101001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01110010101001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01110010101001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01110010101001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01110010101001101011) && ({row_reg, col_reg}<20'b01110010110100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01110010110100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01110010110100011111) && ({row_reg, col_reg}<20'b01110010110101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01110010110101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01110010110101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01110010110101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01110010110101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01110010110101010000) && ({row_reg, col_reg}<20'b01110010111000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01110010111000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01110010111000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01110010111000111000) && ({row_reg, col_reg}<20'b01110010111000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01110010111000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01110010111000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01110010111000111100) && ({row_reg, col_reg}<20'b01110010111000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01110010111000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01110010111000111111) && ({row_reg, col_reg}<20'b01110010111001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01110010111001100110) && ({row_reg, col_reg}<20'b01110010111001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01110010111001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01110010111001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01110010111001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01110010111001101011) && ({row_reg, col_reg}<20'b01110011000100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01110011000100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01110011000100011111) && ({row_reg, col_reg}<20'b01110011000101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01110011000101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01110011000101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01110011000101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01110011000101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01110011000101010000) && ({row_reg, col_reg}<20'b01110011001000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01110011001000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01110011001000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01110011001000111000) && ({row_reg, col_reg}<20'b01110011001000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01110011001000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01110011001000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01110011001000111100) && ({row_reg, col_reg}<20'b01110011001000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01110011001000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01110011001000111111) && ({row_reg, col_reg}<20'b01110011001001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01110011001001100110) && ({row_reg, col_reg}<20'b01110011001001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01110011001001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01110011001001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01110011001001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01110011001001101011) && ({row_reg, col_reg}<20'b01110011010100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01110011010100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01110011010100011111) && ({row_reg, col_reg}<20'b01110011010101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01110011010101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01110011010101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01110011010101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01110011010101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01110011010101010000) && ({row_reg, col_reg}<20'b01110011011000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01110011011000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01110011011000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01110011011000111000) && ({row_reg, col_reg}<20'b01110011011000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01110011011000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01110011011000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01110011011000111100) && ({row_reg, col_reg}<20'b01110011011000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01110011011000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01110011011000111111) && ({row_reg, col_reg}<20'b01110011011001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01110011011001100110) && ({row_reg, col_reg}<20'b01110011011001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01110011011001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01110011011001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01110011011001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01110011011001101011) && ({row_reg, col_reg}<20'b01110011100100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01110011100100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01110011100100011111) && ({row_reg, col_reg}<20'b01110011100101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01110011100101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01110011100101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01110011100101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01110011100101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01110011100101010000) && ({row_reg, col_reg}<20'b01110011101000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01110011101000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01110011101000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01110011101000111000) && ({row_reg, col_reg}<20'b01110011101000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01110011101000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01110011101000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01110011101000111100) && ({row_reg, col_reg}<20'b01110011101000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01110011101000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01110011101000111111) && ({row_reg, col_reg}<20'b01110011101001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01110011101001100110) && ({row_reg, col_reg}<20'b01110011101001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01110011101001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01110011101001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01110011101001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01110011101001101011) && ({row_reg, col_reg}<20'b01110011110100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01110011110100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01110011110100011111) && ({row_reg, col_reg}<20'b01110011110101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01110011110101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01110011110101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01110011110101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01110011110101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01110011110101010000) && ({row_reg, col_reg}<20'b01110011111000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01110011111000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01110011111000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01110011111000111000) && ({row_reg, col_reg}<20'b01110011111000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01110011111000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01110011111000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01110011111000111100) && ({row_reg, col_reg}<20'b01110011111000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01110011111000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01110011111000111111) && ({row_reg, col_reg}<20'b01110011111001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01110011111001100110) && ({row_reg, col_reg}<20'b01110011111001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01110011111001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01110011111001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01110011111001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01110011111001101011) && ({row_reg, col_reg}<20'b01110100000100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01110100000100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01110100000100011111) && ({row_reg, col_reg}<20'b01110100000101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01110100000101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01110100000101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01110100000101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01110100000101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01110100000101010000) && ({row_reg, col_reg}<20'b01110100001000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01110100001000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01110100001000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01110100001000111000) && ({row_reg, col_reg}<20'b01110100001000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01110100001000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01110100001000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01110100001000111100) && ({row_reg, col_reg}<20'b01110100001000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01110100001000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01110100001000111111) && ({row_reg, col_reg}<20'b01110100001001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01110100001001100110) && ({row_reg, col_reg}<20'b01110100001001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01110100001001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01110100001001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01110100001001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01110100001001101011) && ({row_reg, col_reg}<20'b01110100010100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01110100010100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01110100010100011111) && ({row_reg, col_reg}<20'b01110100010101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01110100010101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01110100010101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01110100010101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01110100010101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01110100010101010000) && ({row_reg, col_reg}<20'b01110100011000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01110100011000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01110100011000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01110100011000111000) && ({row_reg, col_reg}<20'b01110100011000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01110100011000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01110100011000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01110100011000111100) && ({row_reg, col_reg}<20'b01110100011000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01110100011000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01110100011000111111) && ({row_reg, col_reg}<20'b01110100011001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01110100011001100110) && ({row_reg, col_reg}<20'b01110100011001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01110100011001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01110100011001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01110100011001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01110100011001101011) && ({row_reg, col_reg}<20'b01110100100100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01110100100100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01110100100100011111) && ({row_reg, col_reg}<20'b01110100100101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01110100100101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01110100100101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01110100100101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01110100100101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01110100100101010000) && ({row_reg, col_reg}<20'b01110100101000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01110100101000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01110100101000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01110100101000111000) && ({row_reg, col_reg}<20'b01110100101000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01110100101000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01110100101000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01110100101000111100) && ({row_reg, col_reg}<20'b01110100101000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01110100101000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01110100101000111111) && ({row_reg, col_reg}<20'b01110100101001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01110100101001100110) && ({row_reg, col_reg}<20'b01110100101001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01110100101001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01110100101001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01110100101001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01110100101001101011) && ({row_reg, col_reg}<20'b01110100110100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01110100110100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01110100110100011111) && ({row_reg, col_reg}<20'b01110100110101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01110100110101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01110100110101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01110100110101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01110100110101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01110100110101010000) && ({row_reg, col_reg}<20'b01110100111000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01110100111000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01110100111000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01110100111000111000) && ({row_reg, col_reg}<20'b01110100111000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01110100111000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01110100111000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01110100111000111100) && ({row_reg, col_reg}<20'b01110100111000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01110100111000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01110100111000111111) && ({row_reg, col_reg}<20'b01110100111001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01110100111001100110) && ({row_reg, col_reg}<20'b01110100111001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01110100111001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01110100111001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01110100111001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01110100111001101011) && ({row_reg, col_reg}<20'b01110101000100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01110101000100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01110101000100011111) && ({row_reg, col_reg}<20'b01110101000101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01110101000101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01110101000101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01110101000101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01110101000101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01110101000101010000) && ({row_reg, col_reg}<20'b01110101001000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01110101001000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01110101001000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01110101001000111000) && ({row_reg, col_reg}<20'b01110101001000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01110101001000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01110101001000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01110101001000111100) && ({row_reg, col_reg}<20'b01110101001000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01110101001000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01110101001000111111) && ({row_reg, col_reg}<20'b01110101001001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01110101001001100110) && ({row_reg, col_reg}<20'b01110101001001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01110101001001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01110101001001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01110101001001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01110101001001101011) && ({row_reg, col_reg}<20'b01110101010100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01110101010100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01110101010100011111) && ({row_reg, col_reg}<20'b01110101010101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01110101010101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01110101010101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01110101010101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01110101010101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01110101010101010000) && ({row_reg, col_reg}<20'b01110101011000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01110101011000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01110101011000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01110101011000111000) && ({row_reg, col_reg}<20'b01110101011000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01110101011000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01110101011000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01110101011000111100) && ({row_reg, col_reg}<20'b01110101011000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01110101011000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01110101011000111111) && ({row_reg, col_reg}<20'b01110101011001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01110101011001100110) && ({row_reg, col_reg}<20'b01110101011001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01110101011001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01110101011001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01110101011001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01110101011001101011) && ({row_reg, col_reg}<20'b01110101100100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01110101100100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01110101100100011111) && ({row_reg, col_reg}<20'b01110101100101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01110101100101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01110101100101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01110101100101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01110101100101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01110101100101010000) && ({row_reg, col_reg}<20'b01110101101000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01110101101000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01110101101000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01110101101000111000) && ({row_reg, col_reg}<20'b01110101101000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01110101101000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01110101101000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01110101101000111100) && ({row_reg, col_reg}<20'b01110101101000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01110101101000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01110101101000111111) && ({row_reg, col_reg}<20'b01110101101001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01110101101001100110) && ({row_reg, col_reg}<20'b01110101101001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01110101101001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01110101101001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01110101101001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01110101101001101011) && ({row_reg, col_reg}<20'b01110101110100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01110101110100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01110101110100011111) && ({row_reg, col_reg}<20'b01110101110101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01110101110101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01110101110101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01110101110101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01110101110101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01110101110101010000) && ({row_reg, col_reg}<20'b01110101111000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01110101111000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01110101111000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01110101111000111000) && ({row_reg, col_reg}<20'b01110101111000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01110101111000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01110101111000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01110101111000111100) && ({row_reg, col_reg}<20'b01110101111000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01110101111000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01110101111000111111) && ({row_reg, col_reg}<20'b01110101111001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01110101111001100110) && ({row_reg, col_reg}<20'b01110101111001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01110101111001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01110101111001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01110101111001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01110101111001101011) && ({row_reg, col_reg}<20'b01110110000100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01110110000100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01110110000100011111) && ({row_reg, col_reg}<20'b01110110000101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01110110000101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01110110000101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01110110000101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01110110000101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01110110000101010000) && ({row_reg, col_reg}<20'b01110110001000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01110110001000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01110110001000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01110110001000111000) && ({row_reg, col_reg}<20'b01110110001000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01110110001000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01110110001000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01110110001000111100) && ({row_reg, col_reg}<20'b01110110001000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01110110001000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01110110001000111111) && ({row_reg, col_reg}<20'b01110110001001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01110110001001100110) && ({row_reg, col_reg}<20'b01110110001001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01110110001001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01110110001001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01110110001001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01110110001001101011) && ({row_reg, col_reg}<20'b01110110010100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01110110010100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01110110010100011111) && ({row_reg, col_reg}<20'b01110110010101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01110110010101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01110110010101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01110110010101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01110110010101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01110110010101010000) && ({row_reg, col_reg}<20'b01110110011000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01110110011000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01110110011000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01110110011000111000) && ({row_reg, col_reg}<20'b01110110011000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01110110011000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01110110011000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01110110011000111100) && ({row_reg, col_reg}<20'b01110110011000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01110110011000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01110110011000111111) && ({row_reg, col_reg}<20'b01110110011001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01110110011001100110) && ({row_reg, col_reg}<20'b01110110011001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01110110011001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01110110011001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01110110011001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01110110011001101011) && ({row_reg, col_reg}<20'b01110110100100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01110110100100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01110110100100011111) && ({row_reg, col_reg}<20'b01110110100101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01110110100101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01110110100101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01110110100101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01110110100101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01110110100101010000) && ({row_reg, col_reg}<20'b01110110101000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01110110101000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01110110101000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01110110101000111000) && ({row_reg, col_reg}<20'b01110110101000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01110110101000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01110110101000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01110110101000111100) && ({row_reg, col_reg}<20'b01110110101000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01110110101000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01110110101000111111) && ({row_reg, col_reg}<20'b01110110101001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01110110101001100110) && ({row_reg, col_reg}<20'b01110110101001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01110110101001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01110110101001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01110110101001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01110110101001101011) && ({row_reg, col_reg}<20'b01110110110100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01110110110100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01110110110100011111) && ({row_reg, col_reg}<20'b01110110110101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01110110110101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01110110110101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01110110110101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01110110110101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01110110110101010000) && ({row_reg, col_reg}<20'b01110110111000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01110110111000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01110110111000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01110110111000111000) && ({row_reg, col_reg}<20'b01110110111000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01110110111000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01110110111000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01110110111000111100) && ({row_reg, col_reg}<20'b01110110111000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01110110111000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01110110111000111111) && ({row_reg, col_reg}<20'b01110110111001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01110110111001100110) && ({row_reg, col_reg}<20'b01110110111001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01110110111001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01110110111001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01110110111001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01110110111001101011) && ({row_reg, col_reg}<20'b01110111000100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01110111000100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01110111000100011111) && ({row_reg, col_reg}<20'b01110111000101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01110111000101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01110111000101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01110111000101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01110111000101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01110111000101010000) && ({row_reg, col_reg}<20'b01110111001000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01110111001000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01110111001000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01110111001000111000) && ({row_reg, col_reg}<20'b01110111001000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01110111001000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01110111001000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01110111001000111100) && ({row_reg, col_reg}<20'b01110111001000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01110111001000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01110111001000111111) && ({row_reg, col_reg}<20'b01110111001001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01110111001001100110) && ({row_reg, col_reg}<20'b01110111001001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01110111001001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01110111001001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01110111001001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01110111001001101011) && ({row_reg, col_reg}<20'b01110111010100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01110111010100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01110111010100011111) && ({row_reg, col_reg}<20'b01110111010101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01110111010101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01110111010101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01110111010101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01110111010101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01110111010101010000) && ({row_reg, col_reg}<20'b01110111011000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01110111011000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01110111011000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01110111011000111000) && ({row_reg, col_reg}<20'b01110111011000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01110111011000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01110111011000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01110111011000111100) && ({row_reg, col_reg}<20'b01110111011000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01110111011000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01110111011000111111) && ({row_reg, col_reg}<20'b01110111011001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01110111011001100110) && ({row_reg, col_reg}<20'b01110111011001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01110111011001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01110111011001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01110111011001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01110111011001101011) && ({row_reg, col_reg}<20'b01110111100100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01110111100100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01110111100100011111) && ({row_reg, col_reg}<20'b01110111100101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01110111100101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01110111100101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01110111100101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01110111100101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01110111100101010000) && ({row_reg, col_reg}<20'b01110111101000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01110111101000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01110111101000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01110111101000111000) && ({row_reg, col_reg}<20'b01110111101000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01110111101000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01110111101000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01110111101000111100) && ({row_reg, col_reg}<20'b01110111101000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01110111101000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01110111101000111111) && ({row_reg, col_reg}<20'b01110111101001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01110111101001100110) && ({row_reg, col_reg}<20'b01110111101001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01110111101001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01110111101001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01110111101001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01110111101001101011) && ({row_reg, col_reg}<20'b01110111110100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01110111110100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01110111110100011111) && ({row_reg, col_reg}<20'b01110111110101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01110111110101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01110111110101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01110111110101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01110111110101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01110111110101010000) && ({row_reg, col_reg}<20'b01110111111000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01110111111000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01110111111000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01110111111000111000) && ({row_reg, col_reg}<20'b01110111111000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01110111111000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01110111111000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01110111111000111100) && ({row_reg, col_reg}<20'b01110111111000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01110111111000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01110111111000111111) && ({row_reg, col_reg}<20'b01110111111001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01110111111001100110) && ({row_reg, col_reg}<20'b01110111111001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01110111111001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01110111111001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01110111111001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01110111111001101011) && ({row_reg, col_reg}<20'b01111000000100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01111000000100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01111000000100011111) && ({row_reg, col_reg}<20'b01111000000101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01111000000101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01111000000101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01111000000101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01111000000101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01111000000101010000) && ({row_reg, col_reg}<20'b01111000001000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01111000001000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01111000001000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01111000001000111000) && ({row_reg, col_reg}<20'b01111000001000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01111000001000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01111000001000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01111000001000111100) && ({row_reg, col_reg}<20'b01111000001000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01111000001000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01111000001000111111) && ({row_reg, col_reg}<20'b01111000001001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01111000001001100110) && ({row_reg, col_reg}<20'b01111000001001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01111000001001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01111000001001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01111000001001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01111000001001101011) && ({row_reg, col_reg}<20'b01111000010100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01111000010100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01111000010100011111) && ({row_reg, col_reg}<20'b01111000010101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01111000010101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01111000010101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01111000010101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01111000010101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01111000010101010000) && ({row_reg, col_reg}<20'b01111000011000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01111000011000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01111000011000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01111000011000111000) && ({row_reg, col_reg}<20'b01111000011000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01111000011000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01111000011000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01111000011000111100) && ({row_reg, col_reg}<20'b01111000011000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01111000011000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01111000011000111111) && ({row_reg, col_reg}<20'b01111000011001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01111000011001100110) && ({row_reg, col_reg}<20'b01111000011001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01111000011001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01111000011001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01111000011001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01111000011001101011) && ({row_reg, col_reg}<20'b01111000100100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01111000100100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01111000100100011111) && ({row_reg, col_reg}<20'b01111000100101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01111000100101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01111000100101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01111000100101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01111000100101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01111000100101010000) && ({row_reg, col_reg}<20'b01111000101000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01111000101000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01111000101000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01111000101000111000) && ({row_reg, col_reg}<20'b01111000101000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01111000101000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01111000101000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01111000101000111100) && ({row_reg, col_reg}<20'b01111000101000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01111000101000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01111000101000111111) && ({row_reg, col_reg}<20'b01111000101001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01111000101001100110) && ({row_reg, col_reg}<20'b01111000101001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01111000101001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01111000101001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01111000101001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01111000101001101011) && ({row_reg, col_reg}<20'b01111000110100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01111000110100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01111000110100011111) && ({row_reg, col_reg}<20'b01111000110101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01111000110101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01111000110101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01111000110101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01111000110101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01111000110101010000) && ({row_reg, col_reg}<20'b01111000111000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01111000111000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01111000111000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01111000111000111000) && ({row_reg, col_reg}<20'b01111000111000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01111000111000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01111000111000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01111000111000111100) && ({row_reg, col_reg}<20'b01111000111000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01111000111000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01111000111000111111) && ({row_reg, col_reg}<20'b01111000111001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01111000111001100110) && ({row_reg, col_reg}<20'b01111000111001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01111000111001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01111000111001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01111000111001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01111000111001101011) && ({row_reg, col_reg}<20'b01111001000100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01111001000100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01111001000100011111) && ({row_reg, col_reg}<20'b01111001000101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01111001000101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01111001000101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01111001000101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01111001000101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01111001000101010000) && ({row_reg, col_reg}<20'b01111001001000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01111001001000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01111001001000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01111001001000111000) && ({row_reg, col_reg}<20'b01111001001000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01111001001000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01111001001000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01111001001000111100) && ({row_reg, col_reg}<20'b01111001001000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01111001001000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01111001001000111111) && ({row_reg, col_reg}<20'b01111001001001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01111001001001100110) && ({row_reg, col_reg}<20'b01111001001001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01111001001001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01111001001001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01111001001001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01111001001001101011) && ({row_reg, col_reg}<20'b01111001010100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01111001010100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01111001010100011111) && ({row_reg, col_reg}<20'b01111001010101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01111001010101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01111001010101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01111001010101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01111001010101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01111001010101010000) && ({row_reg, col_reg}<20'b01111001011000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01111001011000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01111001011000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01111001011000111000) && ({row_reg, col_reg}<20'b01111001011000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01111001011000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01111001011000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01111001011000111100) && ({row_reg, col_reg}<20'b01111001011000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01111001011000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01111001011000111111) && ({row_reg, col_reg}<20'b01111001011001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01111001011001100110) && ({row_reg, col_reg}<20'b01111001011001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01111001011001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01111001011001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01111001011001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01111001011001101011) && ({row_reg, col_reg}<20'b01111001100100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01111001100100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01111001100100011111) && ({row_reg, col_reg}<20'b01111001100101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01111001100101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01111001100101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01111001100101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01111001100101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01111001100101010000) && ({row_reg, col_reg}<20'b01111001101000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01111001101000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01111001101000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01111001101000111000) && ({row_reg, col_reg}<20'b01111001101000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01111001101000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01111001101000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01111001101000111100) && ({row_reg, col_reg}<20'b01111001101000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01111001101000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01111001101000111111) && ({row_reg, col_reg}<20'b01111001101001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01111001101001100110) && ({row_reg, col_reg}<20'b01111001101001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01111001101001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01111001101001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01111001101001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01111001101001101011) && ({row_reg, col_reg}<20'b01111001110100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01111001110100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01111001110100011111) && ({row_reg, col_reg}<20'b01111001110101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01111001110101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01111001110101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01111001110101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01111001110101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01111001110101010000) && ({row_reg, col_reg}<20'b01111001111000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01111001111000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01111001111000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01111001111000111000) && ({row_reg, col_reg}<20'b01111001111000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01111001111000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01111001111000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01111001111000111100) && ({row_reg, col_reg}<20'b01111001111000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01111001111000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01111001111000111111) && ({row_reg, col_reg}<20'b01111001111001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01111001111001100110) && ({row_reg, col_reg}<20'b01111001111001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01111001111001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01111001111001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01111001111001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01111001111001101011) && ({row_reg, col_reg}<20'b01111010000100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01111010000100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01111010000100011111) && ({row_reg, col_reg}<20'b01111010000101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01111010000101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01111010000101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01111010000101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01111010000101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01111010000101010000) && ({row_reg, col_reg}<20'b01111010001000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01111010001000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01111010001000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01111010001000111000) && ({row_reg, col_reg}<20'b01111010001000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01111010001000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01111010001000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01111010001000111100) && ({row_reg, col_reg}<20'b01111010001000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01111010001000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01111010001000111111) && ({row_reg, col_reg}<20'b01111010001001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01111010001001100110) && ({row_reg, col_reg}<20'b01111010001001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01111010001001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01111010001001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01111010001001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01111010001001101011) && ({row_reg, col_reg}<20'b01111010010100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01111010010100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01111010010100011111) && ({row_reg, col_reg}<20'b01111010010101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01111010010101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01111010010101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01111010010101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01111010010101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01111010010101010000) && ({row_reg, col_reg}<20'b01111010011000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01111010011000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01111010011000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01111010011000111000) && ({row_reg, col_reg}<20'b01111010011000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01111010011000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01111010011000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01111010011000111100) && ({row_reg, col_reg}<20'b01111010011000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01111010011000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01111010011000111111) && ({row_reg, col_reg}<20'b01111010011001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01111010011001100110) && ({row_reg, col_reg}<20'b01111010011001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01111010011001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01111010011001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01111010011001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01111010011001101011) && ({row_reg, col_reg}<20'b01111010100100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01111010100100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01111010100100011111) && ({row_reg, col_reg}<20'b01111010100101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01111010100101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01111010100101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01111010100101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01111010100101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01111010100101010000) && ({row_reg, col_reg}<20'b01111010101000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01111010101000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01111010101000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01111010101000111000) && ({row_reg, col_reg}<20'b01111010101000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01111010101000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01111010101000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01111010101000111100) && ({row_reg, col_reg}<20'b01111010101000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01111010101000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01111010101000111111) && ({row_reg, col_reg}<20'b01111010101001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01111010101001100110) && ({row_reg, col_reg}<20'b01111010101001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01111010101001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01111010101001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01111010101001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01111010101001101011) && ({row_reg, col_reg}<20'b01111010110100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01111010110100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01111010110100011111) && ({row_reg, col_reg}<20'b01111010110101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01111010110101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01111010110101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01111010110101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01111010110101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01111010110101010000) && ({row_reg, col_reg}<20'b01111010111000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01111010111000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01111010111000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01111010111000111000) && ({row_reg, col_reg}<20'b01111010111000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01111010111000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01111010111000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01111010111000111100) && ({row_reg, col_reg}<20'b01111010111000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01111010111000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01111010111000111111) && ({row_reg, col_reg}<20'b01111010111001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01111010111001100110) && ({row_reg, col_reg}<20'b01111010111001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01111010111001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01111010111001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01111010111001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01111010111001101011) && ({row_reg, col_reg}<20'b01111011000100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01111011000100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01111011000100011111) && ({row_reg, col_reg}<20'b01111011000101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01111011000101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01111011000101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01111011000101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01111011000101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01111011000101010000) && ({row_reg, col_reg}<20'b01111011001000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01111011001000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01111011001000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01111011001000111000) && ({row_reg, col_reg}<20'b01111011001000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01111011001000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01111011001000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01111011001000111100) && ({row_reg, col_reg}<20'b01111011001000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01111011001000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01111011001000111111) && ({row_reg, col_reg}<20'b01111011001001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01111011001001100110) && ({row_reg, col_reg}<20'b01111011001001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01111011001001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01111011001001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01111011001001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01111011001001101011) && ({row_reg, col_reg}<20'b01111011010100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01111011010100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01111011010100011111) && ({row_reg, col_reg}<20'b01111011010101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01111011010101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01111011010101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01111011010101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01111011010101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01111011010101010000) && ({row_reg, col_reg}<20'b01111011011000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01111011011000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01111011011000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01111011011000111000) && ({row_reg, col_reg}<20'b01111011011000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01111011011000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01111011011000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01111011011000111100) && ({row_reg, col_reg}<20'b01111011011000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01111011011000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01111011011000111111) && ({row_reg, col_reg}<20'b01111011011001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01111011011001100110) && ({row_reg, col_reg}<20'b01111011011001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01111011011001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01111011011001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01111011011001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01111011011001101011) && ({row_reg, col_reg}<20'b01111011100100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01111011100100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01111011100100011111) && ({row_reg, col_reg}<20'b01111011100101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01111011100101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01111011100101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01111011100101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01111011100101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01111011100101010000) && ({row_reg, col_reg}<20'b01111011101000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01111011101000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01111011101000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01111011101000111000) && ({row_reg, col_reg}<20'b01111011101000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01111011101000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01111011101000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01111011101000111100) && ({row_reg, col_reg}<20'b01111011101000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01111011101000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01111011101000111111) && ({row_reg, col_reg}<20'b01111011101001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01111011101001100110) && ({row_reg, col_reg}<20'b01111011101001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01111011101001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01111011101001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01111011101001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01111011101001101011) && ({row_reg, col_reg}<20'b01111011110100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01111011110100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01111011110100011111) && ({row_reg, col_reg}<20'b01111011110101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01111011110101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01111011110101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01111011110101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01111011110101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01111011110101010000) && ({row_reg, col_reg}<20'b01111011111000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01111011111000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01111011111000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01111011111000111000) && ({row_reg, col_reg}<20'b01111011111000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01111011111000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01111011111000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01111011111000111100) && ({row_reg, col_reg}<20'b01111011111000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01111011111000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01111011111000111111) && ({row_reg, col_reg}<20'b01111011111001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01111011111001100110) && ({row_reg, col_reg}<20'b01111011111001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01111011111001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01111011111001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01111011111001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01111011111001101011) && ({row_reg, col_reg}<20'b01111100000100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01111100000100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01111100000100011111) && ({row_reg, col_reg}<20'b01111100000101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01111100000101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01111100000101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01111100000101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01111100000101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01111100000101010000) && ({row_reg, col_reg}<20'b01111100001000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01111100001000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01111100001000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01111100001000111000) && ({row_reg, col_reg}<20'b01111100001000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01111100001000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01111100001000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01111100001000111100) && ({row_reg, col_reg}<20'b01111100001000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01111100001000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01111100001000111111) && ({row_reg, col_reg}<20'b01111100001001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01111100001001100110) && ({row_reg, col_reg}<20'b01111100001001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01111100001001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01111100001001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01111100001001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01111100001001101011) && ({row_reg, col_reg}<20'b01111100010100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01111100010100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01111100010100011111) && ({row_reg, col_reg}<20'b01111100010101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01111100010101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01111100010101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01111100010101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01111100010101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01111100010101010000) && ({row_reg, col_reg}<20'b01111100011000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01111100011000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01111100011000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01111100011000111000) && ({row_reg, col_reg}<20'b01111100011000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01111100011000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01111100011000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01111100011000111100) && ({row_reg, col_reg}<20'b01111100011000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01111100011000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01111100011000111111) && ({row_reg, col_reg}<20'b01111100011001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01111100011001100110) && ({row_reg, col_reg}<20'b01111100011001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01111100011001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01111100011001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01111100011001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01111100011001101011) && ({row_reg, col_reg}<20'b01111100100100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01111100100100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01111100100100011111) && ({row_reg, col_reg}<20'b01111100100101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01111100100101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01111100100101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01111100100101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01111100100101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01111100100101010000) && ({row_reg, col_reg}<20'b01111100101000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01111100101000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01111100101000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01111100101000111000) && ({row_reg, col_reg}<20'b01111100101000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01111100101000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01111100101000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01111100101000111100) && ({row_reg, col_reg}<20'b01111100101000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01111100101000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01111100101000111111) && ({row_reg, col_reg}<20'b01111100101001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01111100101001100110) && ({row_reg, col_reg}<20'b01111100101001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01111100101001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01111100101001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01111100101001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01111100101001101011) && ({row_reg, col_reg}<20'b01111100110100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01111100110100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01111100110100011111) && ({row_reg, col_reg}<20'b01111100110101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01111100110101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01111100110101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01111100110101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01111100110101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01111100110101010000) && ({row_reg, col_reg}<20'b01111100111000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01111100111000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01111100111000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01111100111000111000) && ({row_reg, col_reg}<20'b01111100111000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01111100111000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01111100111000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01111100111000111100) && ({row_reg, col_reg}<20'b01111100111000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01111100111000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01111100111000111111) && ({row_reg, col_reg}<20'b01111100111001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01111100111001100110) && ({row_reg, col_reg}<20'b01111100111001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01111100111001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01111100111001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01111100111001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01111100111001101011) && ({row_reg, col_reg}<20'b01111101000100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01111101000100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01111101000100011111) && ({row_reg, col_reg}<20'b01111101000101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01111101000101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01111101000101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01111101000101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01111101000101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01111101000101010000) && ({row_reg, col_reg}<20'b01111101001000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01111101001000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01111101001000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01111101001000111000) && ({row_reg, col_reg}<20'b01111101001000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01111101001000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01111101001000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01111101001000111100) && ({row_reg, col_reg}<20'b01111101001000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01111101001000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01111101001000111111) && ({row_reg, col_reg}<20'b01111101001001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01111101001001100110) && ({row_reg, col_reg}<20'b01111101001001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01111101001001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01111101001001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01111101001001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01111101001001101011) && ({row_reg, col_reg}<20'b01111101010100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01111101010100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01111101010100011111) && ({row_reg, col_reg}<20'b01111101010101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01111101010101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01111101010101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01111101010101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01111101010101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01111101010101010000) && ({row_reg, col_reg}<20'b01111101011000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01111101011000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01111101011000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01111101011000111000) && ({row_reg, col_reg}<20'b01111101011000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01111101011000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01111101011000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01111101011000111100) && ({row_reg, col_reg}<20'b01111101011000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01111101011000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01111101011000111111) && ({row_reg, col_reg}<20'b01111101011001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01111101011001100110) && ({row_reg, col_reg}<20'b01111101011001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01111101011001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01111101011001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01111101011001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01111101011001101011) && ({row_reg, col_reg}<20'b01111101100100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01111101100100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01111101100100011111) && ({row_reg, col_reg}<20'b01111101100101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01111101100101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01111101100101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01111101100101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01111101100101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01111101100101010000) && ({row_reg, col_reg}<20'b01111101101000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01111101101000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01111101101000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01111101101000111000) && ({row_reg, col_reg}<20'b01111101101000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01111101101000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01111101101000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01111101101000111100) && ({row_reg, col_reg}<20'b01111101101000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01111101101000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01111101101000111111) && ({row_reg, col_reg}<20'b01111101101001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01111101101001100110) && ({row_reg, col_reg}<20'b01111101101001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01111101101001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01111101101001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01111101101001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01111101101001101011) && ({row_reg, col_reg}<20'b01111101110100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01111101110100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01111101110100011111) && ({row_reg, col_reg}<20'b01111101110101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01111101110101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01111101110101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01111101110101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01111101110101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01111101110101010000) && ({row_reg, col_reg}<20'b01111101111000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01111101111000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01111101111000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01111101111000111000) && ({row_reg, col_reg}<20'b01111101111000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01111101111000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01111101111000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01111101111000111100) && ({row_reg, col_reg}<20'b01111101111000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01111101111000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01111101111000111111) && ({row_reg, col_reg}<20'b01111101111001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01111101111001100110) && ({row_reg, col_reg}<20'b01111101111001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01111101111001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01111101111001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01111101111001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01111101111001101011) && ({row_reg, col_reg}<20'b01111110000100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01111110000100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01111110000100011111) && ({row_reg, col_reg}<20'b01111110000101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01111110000101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01111110000101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01111110000101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01111110000101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01111110000101010000) && ({row_reg, col_reg}<20'b01111110001000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01111110001000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01111110001000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01111110001000111000) && ({row_reg, col_reg}<20'b01111110001000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01111110001000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01111110001000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01111110001000111100) && ({row_reg, col_reg}<20'b01111110001000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01111110001000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01111110001000111111) && ({row_reg, col_reg}<20'b01111110001001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01111110001001100110) && ({row_reg, col_reg}<20'b01111110001001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01111110001001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01111110001001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01111110001001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01111110001001101011) && ({row_reg, col_reg}<20'b01111110010100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01111110010100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01111110010100011111) && ({row_reg, col_reg}<20'b01111110010101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01111110010101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01111110010101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01111110010101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01111110010101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01111110010101010000) && ({row_reg, col_reg}<20'b01111110011000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01111110011000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01111110011000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01111110011000111000) && ({row_reg, col_reg}<20'b01111110011000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01111110011000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01111110011000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01111110011000111100) && ({row_reg, col_reg}<20'b01111110011000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01111110011000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01111110011000111111) && ({row_reg, col_reg}<20'b01111110011001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01111110011001100110) && ({row_reg, col_reg}<20'b01111110011001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01111110011001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01111110011001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01111110011001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01111110011001101011) && ({row_reg, col_reg}<20'b01111110100100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01111110100100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01111110100100011111) && ({row_reg, col_reg}<20'b01111110100101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01111110100101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01111110100101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01111110100101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01111110100101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01111110100101010000) && ({row_reg, col_reg}<20'b01111110101000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01111110101000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01111110101000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01111110101000111000) && ({row_reg, col_reg}<20'b01111110101000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01111110101000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01111110101000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01111110101000111100) && ({row_reg, col_reg}<20'b01111110101000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01111110101000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01111110101000111111) && ({row_reg, col_reg}<20'b01111110101001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01111110101001100110) && ({row_reg, col_reg}<20'b01111110101001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01111110101001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01111110101001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01111110101001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01111110101001101011) && ({row_reg, col_reg}<20'b01111110110100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01111110110100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01111110110100011111) && ({row_reg, col_reg}<20'b01111110110101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01111110110101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01111110110101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01111110110101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01111110110101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01111110110101010000) && ({row_reg, col_reg}<20'b01111110111000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01111110111000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01111110111000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01111110111000111000) && ({row_reg, col_reg}<20'b01111110111000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01111110111000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01111110111000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01111110111000111100) && ({row_reg, col_reg}<20'b01111110111000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01111110111000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01111110111000111111) && ({row_reg, col_reg}<20'b01111110111001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01111110111001100110) && ({row_reg, col_reg}<20'b01111110111001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01111110111001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01111110111001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01111110111001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01111110111001101011) && ({row_reg, col_reg}<20'b01111111000100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01111111000100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01111111000100011111) && ({row_reg, col_reg}<20'b01111111000101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01111111000101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01111111000101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01111111000101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01111111000101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01111111000101010000) && ({row_reg, col_reg}<20'b01111111001000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01111111001000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01111111001000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01111111001000111000) && ({row_reg, col_reg}<20'b01111111001000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01111111001000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01111111001000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01111111001000111100) && ({row_reg, col_reg}<20'b01111111001000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01111111001000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01111111001000111111) && ({row_reg, col_reg}<20'b01111111001001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01111111001001100110) && ({row_reg, col_reg}<20'b01111111001001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01111111001001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01111111001001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01111111001001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01111111001001101011) && ({row_reg, col_reg}<20'b01111111010100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01111111010100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01111111010100011111) && ({row_reg, col_reg}<20'b01111111010101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01111111010101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01111111010101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01111111010101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01111111010101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01111111010101010000) && ({row_reg, col_reg}<20'b01111111011000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01111111011000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01111111011000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01111111011000111000) && ({row_reg, col_reg}<20'b01111111011000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01111111011000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01111111011000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01111111011000111100) && ({row_reg, col_reg}<20'b01111111011000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01111111011000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01111111011000111111) && ({row_reg, col_reg}<20'b01111111011001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01111111011001100110) && ({row_reg, col_reg}<20'b01111111011001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01111111011001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01111111011001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01111111011001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01111111011001101011) && ({row_reg, col_reg}<20'b01111111100100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01111111100100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01111111100100011111) && ({row_reg, col_reg}<20'b01111111100101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01111111100101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01111111100101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01111111100101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01111111100101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01111111100101010000) && ({row_reg, col_reg}<20'b01111111101000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01111111101000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01111111101000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01111111101000111000) && ({row_reg, col_reg}<20'b01111111101000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01111111101000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01111111101000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01111111101000111100) && ({row_reg, col_reg}<20'b01111111101000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01111111101000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01111111101000111111) && ({row_reg, col_reg}<20'b01111111101001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01111111101001100110) && ({row_reg, col_reg}<20'b01111111101001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01111111101001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01111111101001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01111111101001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01111111101001101011) && ({row_reg, col_reg}<20'b01111111110100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01111111110100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b01111111110100011111) && ({row_reg, col_reg}<20'b01111111110101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01111111110101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01111111110101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01111111110101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01111111110101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01111111110101010000) && ({row_reg, col_reg}<20'b01111111111000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01111111111000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b01111111111000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b01111111111000111000) && ({row_reg, col_reg}<20'b01111111111000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01111111111000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01111111111000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01111111111000111100) && ({row_reg, col_reg}<20'b01111111111000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b01111111111000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b01111111111000111111) && ({row_reg, col_reg}<20'b01111111111001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b01111111111001100110) && ({row_reg, col_reg}<20'b01111111111001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b01111111111001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b01111111111001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b01111111111001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b01111111111001101011) && ({row_reg, col_reg}<20'b10000000000100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10000000000100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10000000000100011111) && ({row_reg, col_reg}<20'b10000000000101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10000000000101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10000000000101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10000000000101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10000000000101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10000000000101010000) && ({row_reg, col_reg}<20'b10000000001000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10000000001000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10000000001000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10000000001000111000) && ({row_reg, col_reg}<20'b10000000001000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10000000001000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10000000001000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10000000001000111100) && ({row_reg, col_reg}<20'b10000000001000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10000000001000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10000000001000111111) && ({row_reg, col_reg}<20'b10000000001001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10000000001001100110) && ({row_reg, col_reg}<20'b10000000001001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10000000001001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10000000001001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10000000001001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10000000001001101011) && ({row_reg, col_reg}<20'b10000000010100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10000000010100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10000000010100011111) && ({row_reg, col_reg}<20'b10000000010101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10000000010101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10000000010101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10000000010101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10000000010101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10000000010101010000) && ({row_reg, col_reg}<20'b10000000011000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10000000011000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10000000011000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10000000011000111000) && ({row_reg, col_reg}<20'b10000000011000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10000000011000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10000000011000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10000000011000111100) && ({row_reg, col_reg}<20'b10000000011000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10000000011000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10000000011000111111) && ({row_reg, col_reg}<20'b10000000011001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10000000011001100110) && ({row_reg, col_reg}<20'b10000000011001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10000000011001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10000000011001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10000000011001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10000000011001101011) && ({row_reg, col_reg}<20'b10000000100100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10000000100100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10000000100100011111) && ({row_reg, col_reg}<20'b10000000100101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10000000100101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10000000100101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10000000100101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10000000100101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10000000100101010000) && ({row_reg, col_reg}<20'b10000000101000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10000000101000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10000000101000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10000000101000111000) && ({row_reg, col_reg}<20'b10000000101000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10000000101000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10000000101000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10000000101000111100) && ({row_reg, col_reg}<20'b10000000101000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10000000101000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10000000101000111111) && ({row_reg, col_reg}<20'b10000000101001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10000000101001100110) && ({row_reg, col_reg}<20'b10000000101001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10000000101001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10000000101001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10000000101001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10000000101001101011) && ({row_reg, col_reg}<20'b10000000110100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10000000110100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10000000110100011111) && ({row_reg, col_reg}<20'b10000000110101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10000000110101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10000000110101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10000000110101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10000000110101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10000000110101010000) && ({row_reg, col_reg}<20'b10000000111000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10000000111000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10000000111000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10000000111000111000) && ({row_reg, col_reg}<20'b10000000111000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10000000111000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10000000111000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10000000111000111100) && ({row_reg, col_reg}<20'b10000000111000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10000000111000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10000000111000111111) && ({row_reg, col_reg}<20'b10000000111001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10000000111001100110) && ({row_reg, col_reg}<20'b10000000111001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10000000111001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10000000111001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10000000111001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10000000111001101011) && ({row_reg, col_reg}<20'b10000001000100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10000001000100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10000001000100011111) && ({row_reg, col_reg}<20'b10000001000101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10000001000101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10000001000101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10000001000101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10000001000101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10000001000101010000) && ({row_reg, col_reg}<20'b10000001001000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10000001001000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10000001001000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10000001001000111000) && ({row_reg, col_reg}<20'b10000001001000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10000001001000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10000001001000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10000001001000111100) && ({row_reg, col_reg}<20'b10000001001000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10000001001000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10000001001000111111) && ({row_reg, col_reg}<20'b10000001001001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10000001001001100110) && ({row_reg, col_reg}<20'b10000001001001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10000001001001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10000001001001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10000001001001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10000001001001101011) && ({row_reg, col_reg}<20'b10000001010100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10000001010100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10000001010100011111) && ({row_reg, col_reg}<20'b10000001010101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10000001010101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10000001010101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10000001010101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10000001010101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10000001010101010000) && ({row_reg, col_reg}<20'b10000001011000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10000001011000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10000001011000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10000001011000111000) && ({row_reg, col_reg}<20'b10000001011000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10000001011000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10000001011000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10000001011000111100) && ({row_reg, col_reg}<20'b10000001011000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10000001011000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10000001011000111111) && ({row_reg, col_reg}<20'b10000001011001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10000001011001100110) && ({row_reg, col_reg}<20'b10000001011001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10000001011001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10000001011001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10000001011001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10000001011001101011) && ({row_reg, col_reg}<20'b10000001100100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10000001100100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10000001100100011111) && ({row_reg, col_reg}<20'b10000001100101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10000001100101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10000001100101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10000001100101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10000001100101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10000001100101010000) && ({row_reg, col_reg}<20'b10000001101000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10000001101000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10000001101000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10000001101000111000) && ({row_reg, col_reg}<20'b10000001101000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10000001101000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10000001101000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10000001101000111100) && ({row_reg, col_reg}<20'b10000001101000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10000001101000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10000001101000111111) && ({row_reg, col_reg}<20'b10000001101001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10000001101001100110) && ({row_reg, col_reg}<20'b10000001101001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10000001101001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10000001101001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10000001101001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10000001101001101011) && ({row_reg, col_reg}<20'b10000001110100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10000001110100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10000001110100011111) && ({row_reg, col_reg}<20'b10000001110101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10000001110101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10000001110101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10000001110101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10000001110101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10000001110101010000) && ({row_reg, col_reg}<20'b10000001111000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10000001111000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10000001111000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10000001111000111000) && ({row_reg, col_reg}<20'b10000001111000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10000001111000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10000001111000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10000001111000111100) && ({row_reg, col_reg}<20'b10000001111000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10000001111000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10000001111000111111) && ({row_reg, col_reg}<20'b10000001111001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10000001111001100110) && ({row_reg, col_reg}<20'b10000001111001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10000001111001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10000001111001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10000001111001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10000001111001101011) && ({row_reg, col_reg}<20'b10000010000100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10000010000100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10000010000100011111) && ({row_reg, col_reg}<20'b10000010000101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10000010000101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10000010000101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10000010000101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10000010000101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10000010000101010000) && ({row_reg, col_reg}<20'b10000010001000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10000010001000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10000010001000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10000010001000111000) && ({row_reg, col_reg}<20'b10000010001000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10000010001000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10000010001000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10000010001000111100) && ({row_reg, col_reg}<20'b10000010001000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10000010001000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10000010001000111111) && ({row_reg, col_reg}<20'b10000010001001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10000010001001100110) && ({row_reg, col_reg}<20'b10000010001001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10000010001001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10000010001001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10000010001001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10000010001001101011) && ({row_reg, col_reg}<20'b10000010010100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10000010010100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10000010010100011111) && ({row_reg, col_reg}<20'b10000010010101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10000010010101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10000010010101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10000010010101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10000010010101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10000010010101010000) && ({row_reg, col_reg}<20'b10000010011000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10000010011000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10000010011000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10000010011000111000) && ({row_reg, col_reg}<20'b10000010011000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10000010011000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10000010011000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10000010011000111100) && ({row_reg, col_reg}<20'b10000010011000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10000010011000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10000010011000111111) && ({row_reg, col_reg}<20'b10000010011001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10000010011001100110) && ({row_reg, col_reg}<20'b10000010011001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10000010011001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10000010011001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10000010011001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10000010011001101011) && ({row_reg, col_reg}<20'b10000010100100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10000010100100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10000010100100011111) && ({row_reg, col_reg}<20'b10000010100101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10000010100101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10000010100101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10000010100101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10000010100101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10000010100101010000) && ({row_reg, col_reg}<20'b10000010101000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10000010101000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10000010101000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10000010101000111000) && ({row_reg, col_reg}<20'b10000010101000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10000010101000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10000010101000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10000010101000111100) && ({row_reg, col_reg}<20'b10000010101000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10000010101000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10000010101000111111) && ({row_reg, col_reg}<20'b10000010101001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10000010101001100110) && ({row_reg, col_reg}<20'b10000010101001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10000010101001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10000010101001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10000010101001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10000010101001101011) && ({row_reg, col_reg}<20'b10000010110100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10000010110100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10000010110100011111) && ({row_reg, col_reg}<20'b10000010110101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10000010110101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10000010110101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10000010110101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10000010110101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10000010110101010000) && ({row_reg, col_reg}<20'b10000010111000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10000010111000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10000010111000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10000010111000111000) && ({row_reg, col_reg}<20'b10000010111000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10000010111000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10000010111000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10000010111000111100) && ({row_reg, col_reg}<20'b10000010111000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10000010111000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10000010111000111111) && ({row_reg, col_reg}<20'b10000010111001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10000010111001100110) && ({row_reg, col_reg}<20'b10000010111001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10000010111001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10000010111001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10000010111001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10000010111001101011) && ({row_reg, col_reg}<20'b10000011000100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10000011000100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10000011000100011111) && ({row_reg, col_reg}<20'b10000011000101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10000011000101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10000011000101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10000011000101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10000011000101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10000011000101010000) && ({row_reg, col_reg}<20'b10000011001000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10000011001000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10000011001000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10000011001000111000) && ({row_reg, col_reg}<20'b10000011001000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10000011001000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10000011001000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10000011001000111100) && ({row_reg, col_reg}<20'b10000011001000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10000011001000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10000011001000111111) && ({row_reg, col_reg}<20'b10000011001001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10000011001001100110) && ({row_reg, col_reg}<20'b10000011001001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10000011001001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10000011001001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10000011001001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10000011001001101011) && ({row_reg, col_reg}<20'b10000011010100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10000011010100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10000011010100011111) && ({row_reg, col_reg}<20'b10000011010101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10000011010101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10000011010101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10000011010101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10000011010101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10000011010101010000) && ({row_reg, col_reg}<20'b10000011011000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10000011011000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10000011011000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10000011011000111000) && ({row_reg, col_reg}<20'b10000011011000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10000011011000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10000011011000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10000011011000111100) && ({row_reg, col_reg}<20'b10000011011000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10000011011000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10000011011000111111) && ({row_reg, col_reg}<20'b10000011011001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10000011011001100110) && ({row_reg, col_reg}<20'b10000011011001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10000011011001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10000011011001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10000011011001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10000011011001101011) && ({row_reg, col_reg}<20'b10000011100100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10000011100100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10000011100100011111) && ({row_reg, col_reg}<20'b10000011100101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10000011100101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10000011100101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10000011100101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10000011100101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10000011100101010000) && ({row_reg, col_reg}<20'b10000011101000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10000011101000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10000011101000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10000011101000111000) && ({row_reg, col_reg}<20'b10000011101000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10000011101000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10000011101000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10000011101000111100) && ({row_reg, col_reg}<20'b10000011101000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10000011101000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10000011101000111111) && ({row_reg, col_reg}<20'b10000011101001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10000011101001100110) && ({row_reg, col_reg}<20'b10000011101001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10000011101001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10000011101001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10000011101001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10000011101001101011) && ({row_reg, col_reg}<20'b10000011110100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10000011110100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10000011110100011111) && ({row_reg, col_reg}<20'b10000011110101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10000011110101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10000011110101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10000011110101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10000011110101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10000011110101010000) && ({row_reg, col_reg}<20'b10000011111000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10000011111000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10000011111000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10000011111000111000) && ({row_reg, col_reg}<20'b10000011111000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10000011111000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10000011111000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10000011111000111100) && ({row_reg, col_reg}<20'b10000011111000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10000011111000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10000011111000111111) && ({row_reg, col_reg}<20'b10000011111001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10000011111001100110) && ({row_reg, col_reg}<20'b10000011111001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10000011111001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10000011111001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10000011111001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10000011111001101011) && ({row_reg, col_reg}<20'b10000100000100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10000100000100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10000100000100011111) && ({row_reg, col_reg}<20'b10000100000101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10000100000101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10000100000101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10000100000101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10000100000101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10000100000101010000) && ({row_reg, col_reg}<20'b10000100001000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10000100001000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10000100001000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10000100001000111000) && ({row_reg, col_reg}<20'b10000100001000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10000100001000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10000100001000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10000100001000111100) && ({row_reg, col_reg}<20'b10000100001000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10000100001000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10000100001000111111) && ({row_reg, col_reg}<20'b10000100001001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10000100001001100110) && ({row_reg, col_reg}<20'b10000100001001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10000100001001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10000100001001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10000100001001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10000100001001101011) && ({row_reg, col_reg}<20'b10000100010100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10000100010100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10000100010100011111) && ({row_reg, col_reg}<20'b10000100010101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10000100010101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10000100010101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10000100010101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10000100010101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10000100010101010000) && ({row_reg, col_reg}<20'b10000100011000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10000100011000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10000100011000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10000100011000111000) && ({row_reg, col_reg}<20'b10000100011000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10000100011000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10000100011000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10000100011000111100) && ({row_reg, col_reg}<20'b10000100011000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10000100011000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10000100011000111111) && ({row_reg, col_reg}<20'b10000100011001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10000100011001100110) && ({row_reg, col_reg}<20'b10000100011001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10000100011001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10000100011001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10000100011001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10000100011001101011) && ({row_reg, col_reg}<20'b10000100100100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10000100100100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10000100100100011111) && ({row_reg, col_reg}<20'b10000100100101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10000100100101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10000100100101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10000100100101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10000100100101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10000100100101010000) && ({row_reg, col_reg}<20'b10000100101000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10000100101000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10000100101000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10000100101000111000) && ({row_reg, col_reg}<20'b10000100101000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10000100101000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10000100101000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10000100101000111100) && ({row_reg, col_reg}<20'b10000100101000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10000100101000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10000100101000111111) && ({row_reg, col_reg}<20'b10000100101001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10000100101001100110) && ({row_reg, col_reg}<20'b10000100101001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10000100101001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10000100101001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10000100101001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10000100101001101011) && ({row_reg, col_reg}<20'b10000100110100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10000100110100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10000100110100011111) && ({row_reg, col_reg}<20'b10000100110101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10000100110101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10000100110101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10000100110101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10000100110101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10000100110101010000) && ({row_reg, col_reg}<20'b10000100111000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10000100111000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10000100111000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10000100111000111000) && ({row_reg, col_reg}<20'b10000100111000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10000100111000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10000100111000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10000100111000111100) && ({row_reg, col_reg}<20'b10000100111000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10000100111000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10000100111000111111) && ({row_reg, col_reg}<20'b10000100111001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10000100111001100110) && ({row_reg, col_reg}<20'b10000100111001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10000100111001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10000100111001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10000100111001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10000100111001101011) && ({row_reg, col_reg}<20'b10000101000100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10000101000100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10000101000100011111) && ({row_reg, col_reg}<20'b10000101000101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10000101000101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10000101000101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10000101000101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10000101000101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10000101000101010000) && ({row_reg, col_reg}<20'b10000101001000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10000101001000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10000101001000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10000101001000111000) && ({row_reg, col_reg}<20'b10000101001000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10000101001000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10000101001000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10000101001000111100) && ({row_reg, col_reg}<20'b10000101001000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10000101001000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10000101001000111111) && ({row_reg, col_reg}<20'b10000101001001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10000101001001100110) && ({row_reg, col_reg}<20'b10000101001001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10000101001001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10000101001001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10000101001001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10000101001001101011) && ({row_reg, col_reg}<20'b10000101010100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10000101010100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10000101010100011111) && ({row_reg, col_reg}<20'b10000101010101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10000101010101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10000101010101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10000101010101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10000101010101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10000101010101010000) && ({row_reg, col_reg}<20'b10000101011000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10000101011000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10000101011000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10000101011000111000) && ({row_reg, col_reg}<20'b10000101011000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10000101011000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10000101011000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10000101011000111100) && ({row_reg, col_reg}<20'b10000101011000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10000101011000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10000101011000111111) && ({row_reg, col_reg}<20'b10000101011001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10000101011001100110) && ({row_reg, col_reg}<20'b10000101011001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10000101011001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10000101011001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10000101011001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10000101011001101011) && ({row_reg, col_reg}<20'b10000101100100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10000101100100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10000101100100011111) && ({row_reg, col_reg}<20'b10000101100101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10000101100101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10000101100101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10000101100101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10000101100101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10000101100101010000) && ({row_reg, col_reg}<20'b10000101101000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10000101101000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10000101101000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10000101101000111000) && ({row_reg, col_reg}<20'b10000101101000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10000101101000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10000101101000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10000101101000111100) && ({row_reg, col_reg}<20'b10000101101000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10000101101000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10000101101000111111) && ({row_reg, col_reg}<20'b10000101101001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10000101101001100110) && ({row_reg, col_reg}<20'b10000101101001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10000101101001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10000101101001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10000101101001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10000101101001101011) && ({row_reg, col_reg}<20'b10000101110100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10000101110100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10000101110100011111) && ({row_reg, col_reg}<20'b10000101110101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10000101110101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10000101110101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10000101110101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10000101110101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10000101110101010000) && ({row_reg, col_reg}<20'b10000101111000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10000101111000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10000101111000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10000101111000111000) && ({row_reg, col_reg}<20'b10000101111000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10000101111000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10000101111000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10000101111000111100) && ({row_reg, col_reg}<20'b10000101111000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10000101111000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10000101111000111111) && ({row_reg, col_reg}<20'b10000101111001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10000101111001100110) && ({row_reg, col_reg}<20'b10000101111001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10000101111001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10000101111001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10000101111001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10000101111001101011) && ({row_reg, col_reg}<20'b10000110000100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10000110000100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10000110000100011111) && ({row_reg, col_reg}<20'b10000110000101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10000110000101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10000110000101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10000110000101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10000110000101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10000110000101010000) && ({row_reg, col_reg}<20'b10000110001000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10000110001000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10000110001000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10000110001000111000) && ({row_reg, col_reg}<20'b10000110001000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10000110001000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10000110001000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10000110001000111100) && ({row_reg, col_reg}<20'b10000110001000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10000110001000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10000110001000111111) && ({row_reg, col_reg}<20'b10000110001001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10000110001001100110) && ({row_reg, col_reg}<20'b10000110001001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10000110001001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10000110001001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10000110001001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10000110001001101011) && ({row_reg, col_reg}<20'b10000110010100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10000110010100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10000110010100011111) && ({row_reg, col_reg}<20'b10000110010101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10000110010101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10000110010101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10000110010101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10000110010101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10000110010101010000) && ({row_reg, col_reg}<20'b10000110011000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10000110011000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10000110011000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10000110011000111000) && ({row_reg, col_reg}<20'b10000110011000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10000110011000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10000110011000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10000110011000111100) && ({row_reg, col_reg}<20'b10000110011000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10000110011000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10000110011000111111) && ({row_reg, col_reg}<20'b10000110011001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10000110011001100110) && ({row_reg, col_reg}<20'b10000110011001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10000110011001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10000110011001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10000110011001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10000110011001101011) && ({row_reg, col_reg}<20'b10000110100100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10000110100100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10000110100100011111) && ({row_reg, col_reg}<20'b10000110100101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10000110100101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10000110100101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10000110100101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10000110100101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10000110100101010000) && ({row_reg, col_reg}<20'b10000110101000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10000110101000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10000110101000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10000110101000111000) && ({row_reg, col_reg}<20'b10000110101000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10000110101000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10000110101000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10000110101000111100) && ({row_reg, col_reg}<20'b10000110101000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10000110101000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10000110101000111111) && ({row_reg, col_reg}<20'b10000110101001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10000110101001100110) && ({row_reg, col_reg}<20'b10000110101001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10000110101001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10000110101001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10000110101001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10000110101001101011) && ({row_reg, col_reg}<20'b10000110110100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10000110110100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10000110110100011111) && ({row_reg, col_reg}<20'b10000110110101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10000110110101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10000110110101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10000110110101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10000110110101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10000110110101010000) && ({row_reg, col_reg}<20'b10000110111000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10000110111000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10000110111000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10000110111000111000) && ({row_reg, col_reg}<20'b10000110111000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10000110111000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10000110111000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10000110111000111100) && ({row_reg, col_reg}<20'b10000110111000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10000110111000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10000110111000111111) && ({row_reg, col_reg}<20'b10000110111001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10000110111001100110) && ({row_reg, col_reg}<20'b10000110111001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10000110111001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10000110111001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10000110111001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10000110111001101011) && ({row_reg, col_reg}<20'b10000111000100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10000111000100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10000111000100011111) && ({row_reg, col_reg}<20'b10000111000101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10000111000101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10000111000101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10000111000101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10000111000101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10000111000101010000) && ({row_reg, col_reg}<20'b10000111001000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10000111001000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10000111001000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10000111001000111000) && ({row_reg, col_reg}<20'b10000111001000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10000111001000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10000111001000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10000111001000111100) && ({row_reg, col_reg}<20'b10000111001000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10000111001000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10000111001000111111) && ({row_reg, col_reg}<20'b10000111001001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10000111001001100110) && ({row_reg, col_reg}<20'b10000111001001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10000111001001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10000111001001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10000111001001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10000111001001101011) && ({row_reg, col_reg}<20'b10000111010100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10000111010100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10000111010100011111) && ({row_reg, col_reg}<20'b10000111010101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10000111010101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10000111010101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10000111010101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10000111010101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10000111010101010000) && ({row_reg, col_reg}<20'b10000111011000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10000111011000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10000111011000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10000111011000111000) && ({row_reg, col_reg}<20'b10000111011000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10000111011000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10000111011000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10000111011000111100) && ({row_reg, col_reg}<20'b10000111011000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10000111011000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10000111011000111111) && ({row_reg, col_reg}<20'b10000111011001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10000111011001100110) && ({row_reg, col_reg}<20'b10000111011001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10000111011001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10000111011001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10000111011001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10000111011001101011) && ({row_reg, col_reg}<20'b10000111100100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10000111100100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10000111100100011111) && ({row_reg, col_reg}<20'b10000111100101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10000111100101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10000111100101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10000111100101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10000111100101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10000111100101010000) && ({row_reg, col_reg}<20'b10000111101000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10000111101000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10000111101000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10000111101000111000) && ({row_reg, col_reg}<20'b10000111101000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10000111101000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10000111101000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10000111101000111100) && ({row_reg, col_reg}<20'b10000111101000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10000111101000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10000111101000111111) && ({row_reg, col_reg}<20'b10000111101001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10000111101001100110) && ({row_reg, col_reg}<20'b10000111101001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10000111101001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10000111101001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10000111101001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10000111101001101011) && ({row_reg, col_reg}<20'b10000111110100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10000111110100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10000111110100011111) && ({row_reg, col_reg}<20'b10000111110101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10000111110101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10000111110101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10000111110101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10000111110101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10000111110101010000) && ({row_reg, col_reg}<20'b10000111111000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10000111111000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10000111111000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10000111111000111000) && ({row_reg, col_reg}<20'b10000111111000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10000111111000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10000111111000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10000111111000111100) && ({row_reg, col_reg}<20'b10000111111000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10000111111000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10000111111000111111) && ({row_reg, col_reg}<20'b10000111111001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10000111111001100110) && ({row_reg, col_reg}<20'b10000111111001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10000111111001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10000111111001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10000111111001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10000111111001101011) && ({row_reg, col_reg}<20'b10001000000100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10001000000100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10001000000100011111) && ({row_reg, col_reg}<20'b10001000000101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10001000000101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10001000000101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10001000000101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10001000000101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10001000000101010000) && ({row_reg, col_reg}<20'b10001000001000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10001000001000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10001000001000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10001000001000111000) && ({row_reg, col_reg}<20'b10001000001000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10001000001000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10001000001000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10001000001000111100) && ({row_reg, col_reg}<20'b10001000001000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10001000001000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10001000001000111111) && ({row_reg, col_reg}<20'b10001000001001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10001000001001100110) && ({row_reg, col_reg}<20'b10001000001001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10001000001001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10001000001001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10001000001001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10001000001001101011) && ({row_reg, col_reg}<20'b10001000010100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10001000010100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10001000010100011111) && ({row_reg, col_reg}<20'b10001000010101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10001000010101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10001000010101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10001000010101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10001000010101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10001000010101010000) && ({row_reg, col_reg}<20'b10001000011000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10001000011000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10001000011000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10001000011000111000) && ({row_reg, col_reg}<20'b10001000011000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10001000011000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10001000011000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10001000011000111100) && ({row_reg, col_reg}<20'b10001000011000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10001000011000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10001000011000111111) && ({row_reg, col_reg}<20'b10001000011001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10001000011001100110) && ({row_reg, col_reg}<20'b10001000011001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10001000011001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10001000011001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10001000011001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10001000011001101011) && ({row_reg, col_reg}<20'b10001000100100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10001000100100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10001000100100011111) && ({row_reg, col_reg}<20'b10001000100101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10001000100101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10001000100101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10001000100101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10001000100101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10001000100101010000) && ({row_reg, col_reg}<20'b10001000101000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10001000101000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10001000101000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10001000101000111000) && ({row_reg, col_reg}<20'b10001000101000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10001000101000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10001000101000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10001000101000111100) && ({row_reg, col_reg}<20'b10001000101000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10001000101000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10001000101000111111) && ({row_reg, col_reg}<20'b10001000101001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10001000101001100110) && ({row_reg, col_reg}<20'b10001000101001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10001000101001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10001000101001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10001000101001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10001000101001101011) && ({row_reg, col_reg}<20'b10001000110100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10001000110100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10001000110100011111) && ({row_reg, col_reg}<20'b10001000110101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10001000110101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10001000110101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10001000110101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10001000110101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10001000110101010000) && ({row_reg, col_reg}<20'b10001000111000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10001000111000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10001000111000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10001000111000111000) && ({row_reg, col_reg}<20'b10001000111000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10001000111000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10001000111000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10001000111000111100) && ({row_reg, col_reg}<20'b10001000111000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10001000111000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10001000111000111111) && ({row_reg, col_reg}<20'b10001000111001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10001000111001100110) && ({row_reg, col_reg}<20'b10001000111001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10001000111001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10001000111001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10001000111001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10001000111001101011) && ({row_reg, col_reg}<20'b10001001000100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10001001000100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10001001000100011111) && ({row_reg, col_reg}<20'b10001001000101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10001001000101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10001001000101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10001001000101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10001001000101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10001001000101010000) && ({row_reg, col_reg}<20'b10001001001000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10001001001000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10001001001000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10001001001000111000) && ({row_reg, col_reg}<20'b10001001001000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10001001001000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10001001001000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10001001001000111100) && ({row_reg, col_reg}<20'b10001001001000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10001001001000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10001001001000111111) && ({row_reg, col_reg}<20'b10001001001001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10001001001001100110) && ({row_reg, col_reg}<20'b10001001001001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10001001001001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10001001001001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10001001001001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10001001001001101011) && ({row_reg, col_reg}<20'b10001001010100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10001001010100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10001001010100011111) && ({row_reg, col_reg}<20'b10001001010101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10001001010101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10001001010101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10001001010101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10001001010101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10001001010101010000) && ({row_reg, col_reg}<20'b10001001011000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10001001011000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10001001011000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10001001011000111000) && ({row_reg, col_reg}<20'b10001001011000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10001001011000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10001001011000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10001001011000111100) && ({row_reg, col_reg}<20'b10001001011000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10001001011000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10001001011000111111) && ({row_reg, col_reg}<20'b10001001011001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10001001011001100110) && ({row_reg, col_reg}<20'b10001001011001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10001001011001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10001001011001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10001001011001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10001001011001101011) && ({row_reg, col_reg}<20'b10001001100100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10001001100100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10001001100100011111) && ({row_reg, col_reg}<20'b10001001100101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10001001100101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10001001100101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10001001100101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10001001100101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10001001100101010000) && ({row_reg, col_reg}<20'b10001001101000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10001001101000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10001001101000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10001001101000111000) && ({row_reg, col_reg}<20'b10001001101000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10001001101000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10001001101000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10001001101000111100) && ({row_reg, col_reg}<20'b10001001101000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10001001101000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10001001101000111111) && ({row_reg, col_reg}<20'b10001001101001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10001001101001100110) && ({row_reg, col_reg}<20'b10001001101001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10001001101001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10001001101001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10001001101001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10001001101001101011) && ({row_reg, col_reg}<20'b10001001110100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10001001110100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10001001110100011111) && ({row_reg, col_reg}<20'b10001001110101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10001001110101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10001001110101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10001001110101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10001001110101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10001001110101010000) && ({row_reg, col_reg}<20'b10001001111000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10001001111000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10001001111000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10001001111000111000) && ({row_reg, col_reg}<20'b10001001111000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10001001111000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10001001111000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10001001111000111100) && ({row_reg, col_reg}<20'b10001001111000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10001001111000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10001001111000111111) && ({row_reg, col_reg}<20'b10001001111001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10001001111001100110) && ({row_reg, col_reg}<20'b10001001111001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10001001111001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10001001111001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10001001111001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10001001111001101011) && ({row_reg, col_reg}<20'b10001010000100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10001010000100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10001010000100011111) && ({row_reg, col_reg}<20'b10001010000101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10001010000101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10001010000101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10001010000101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10001010000101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10001010000101010000) && ({row_reg, col_reg}<20'b10001010001000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10001010001000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10001010001000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10001010001000111000) && ({row_reg, col_reg}<20'b10001010001000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10001010001000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10001010001000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10001010001000111100) && ({row_reg, col_reg}<20'b10001010001000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10001010001000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10001010001000111111) && ({row_reg, col_reg}<20'b10001010001001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10001010001001100110) && ({row_reg, col_reg}<20'b10001010001001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10001010001001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10001010001001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10001010001001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10001010001001101011) && ({row_reg, col_reg}<20'b10001010010100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10001010010100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10001010010100011111) && ({row_reg, col_reg}<20'b10001010010101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10001010010101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10001010010101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10001010010101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10001010010101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10001010010101010000) && ({row_reg, col_reg}<20'b10001010011000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10001010011000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10001010011000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10001010011000111000) && ({row_reg, col_reg}<20'b10001010011000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10001010011000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10001010011000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10001010011000111100) && ({row_reg, col_reg}<20'b10001010011000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10001010011000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10001010011000111111) && ({row_reg, col_reg}<20'b10001010011001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10001010011001100110) && ({row_reg, col_reg}<20'b10001010011001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10001010011001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10001010011001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10001010011001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10001010011001101011) && ({row_reg, col_reg}<20'b10001010100100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10001010100100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10001010100100011111) && ({row_reg, col_reg}<20'b10001010100101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10001010100101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10001010100101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10001010100101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10001010100101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10001010100101010000) && ({row_reg, col_reg}<20'b10001010101000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10001010101000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10001010101000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10001010101000111000) && ({row_reg, col_reg}<20'b10001010101000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10001010101000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10001010101000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10001010101000111100) && ({row_reg, col_reg}<20'b10001010101000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10001010101000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10001010101000111111) && ({row_reg, col_reg}<20'b10001010101001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10001010101001100110) && ({row_reg, col_reg}<20'b10001010101001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10001010101001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10001010101001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10001010101001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10001010101001101011) && ({row_reg, col_reg}<20'b10001010110100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10001010110100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10001010110100011111) && ({row_reg, col_reg}<20'b10001010110101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10001010110101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10001010110101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10001010110101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10001010110101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10001010110101010000) && ({row_reg, col_reg}<20'b10001010111000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10001010111000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10001010111000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10001010111000111000) && ({row_reg, col_reg}<20'b10001010111000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10001010111000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10001010111000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10001010111000111100) && ({row_reg, col_reg}<20'b10001010111000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10001010111000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10001010111000111111) && ({row_reg, col_reg}<20'b10001010111001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10001010111001100110) && ({row_reg, col_reg}<20'b10001010111001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10001010111001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10001010111001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10001010111001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10001010111001101011) && ({row_reg, col_reg}<20'b10001011000100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10001011000100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10001011000100011111) && ({row_reg, col_reg}<20'b10001011000101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10001011000101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10001011000101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10001011000101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10001011000101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10001011000101010000) && ({row_reg, col_reg}<20'b10001011001000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10001011001000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10001011001000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10001011001000111000) && ({row_reg, col_reg}<20'b10001011001000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10001011001000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10001011001000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10001011001000111100) && ({row_reg, col_reg}<20'b10001011001000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10001011001000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10001011001000111111) && ({row_reg, col_reg}<20'b10001011001001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10001011001001100110) && ({row_reg, col_reg}<20'b10001011001001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10001011001001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10001011001001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10001011001001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10001011001001101011) && ({row_reg, col_reg}<20'b10001011010100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10001011010100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10001011010100011111) && ({row_reg, col_reg}<20'b10001011010101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10001011010101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10001011010101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10001011010101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10001011010101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10001011010101010000) && ({row_reg, col_reg}<20'b10001011011000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10001011011000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10001011011000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10001011011000111000) && ({row_reg, col_reg}<20'b10001011011000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10001011011000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10001011011000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10001011011000111100) && ({row_reg, col_reg}<20'b10001011011000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10001011011000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10001011011000111111) && ({row_reg, col_reg}<20'b10001011011001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10001011011001100110) && ({row_reg, col_reg}<20'b10001011011001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10001011011001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10001011011001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10001011011001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10001011011001101011) && ({row_reg, col_reg}<20'b10001011100100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10001011100100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10001011100100011111) && ({row_reg, col_reg}<20'b10001011100101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10001011100101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10001011100101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10001011100101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10001011100101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10001011100101010000) && ({row_reg, col_reg}<20'b10001011101000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10001011101000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10001011101000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10001011101000111000) && ({row_reg, col_reg}<20'b10001011101000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10001011101000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10001011101000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10001011101000111100) && ({row_reg, col_reg}<20'b10001011101000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10001011101000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10001011101000111111) && ({row_reg, col_reg}<20'b10001011101001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10001011101001100110) && ({row_reg, col_reg}<20'b10001011101001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10001011101001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10001011101001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10001011101001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10001011101001101011) && ({row_reg, col_reg}<20'b10001011110100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10001011110100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10001011110100011111) && ({row_reg, col_reg}<20'b10001011110101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10001011110101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10001011110101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10001011110101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10001011110101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10001011110101010000) && ({row_reg, col_reg}<20'b10001011111000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10001011111000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10001011111000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10001011111000111000) && ({row_reg, col_reg}<20'b10001011111000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10001011111000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10001011111000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10001011111000111100) && ({row_reg, col_reg}<20'b10001011111000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10001011111000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10001011111000111111) && ({row_reg, col_reg}<20'b10001011111001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10001011111001100110) && ({row_reg, col_reg}<20'b10001011111001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10001011111001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10001011111001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10001011111001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10001011111001101011) && ({row_reg, col_reg}<20'b10001100000100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10001100000100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10001100000100011111) && ({row_reg, col_reg}<20'b10001100000101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10001100000101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10001100000101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10001100000101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10001100000101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10001100000101010000) && ({row_reg, col_reg}<20'b10001100001000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10001100001000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10001100001000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10001100001000111000) && ({row_reg, col_reg}<20'b10001100001000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10001100001000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10001100001000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10001100001000111100) && ({row_reg, col_reg}<20'b10001100001000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10001100001000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10001100001000111111) && ({row_reg, col_reg}<20'b10001100001001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10001100001001100110) && ({row_reg, col_reg}<20'b10001100001001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10001100001001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10001100001001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10001100001001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10001100001001101011) && ({row_reg, col_reg}<20'b10001100010100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10001100010100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10001100010100011111) && ({row_reg, col_reg}<20'b10001100010101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10001100010101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10001100010101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10001100010101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10001100010101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10001100010101010000) && ({row_reg, col_reg}<20'b10001100011000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10001100011000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10001100011000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10001100011000111000) && ({row_reg, col_reg}<20'b10001100011000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10001100011000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10001100011000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10001100011000111100) && ({row_reg, col_reg}<20'b10001100011000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10001100011000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10001100011000111111) && ({row_reg, col_reg}<20'b10001100011001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10001100011001100110) && ({row_reg, col_reg}<20'b10001100011001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10001100011001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10001100011001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10001100011001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10001100011001101011) && ({row_reg, col_reg}<20'b10001100100100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10001100100100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10001100100100011111) && ({row_reg, col_reg}<20'b10001100100101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10001100100101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10001100100101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10001100100101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10001100100101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10001100100101010000) && ({row_reg, col_reg}<20'b10001100101000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10001100101000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10001100101000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10001100101000111000) && ({row_reg, col_reg}<20'b10001100101000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10001100101000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10001100101000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10001100101000111100) && ({row_reg, col_reg}<20'b10001100101000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10001100101000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10001100101000111111) && ({row_reg, col_reg}<20'b10001100101001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10001100101001100110) && ({row_reg, col_reg}<20'b10001100101001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10001100101001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10001100101001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10001100101001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10001100101001101011) && ({row_reg, col_reg}<20'b10001100110100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10001100110100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10001100110100011111) && ({row_reg, col_reg}<20'b10001100110101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10001100110101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10001100110101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10001100110101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10001100110101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10001100110101010000) && ({row_reg, col_reg}<20'b10001100111000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10001100111000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10001100111000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10001100111000111000) && ({row_reg, col_reg}<20'b10001100111000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10001100111000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10001100111000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10001100111000111100) && ({row_reg, col_reg}<20'b10001100111000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10001100111000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10001100111000111111) && ({row_reg, col_reg}<20'b10001100111001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10001100111001100110) && ({row_reg, col_reg}<20'b10001100111001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10001100111001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10001100111001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10001100111001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10001100111001101011) && ({row_reg, col_reg}<20'b10001101000100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10001101000100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10001101000100011111) && ({row_reg, col_reg}<20'b10001101000101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10001101000101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10001101000101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10001101000101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10001101000101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10001101000101010000) && ({row_reg, col_reg}<20'b10001101001000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10001101001000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10001101001000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10001101001000111000) && ({row_reg, col_reg}<20'b10001101001000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10001101001000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10001101001000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10001101001000111100) && ({row_reg, col_reg}<20'b10001101001000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10001101001000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10001101001000111111) && ({row_reg, col_reg}<20'b10001101001001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10001101001001100110) && ({row_reg, col_reg}<20'b10001101001001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10001101001001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10001101001001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10001101001001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10001101001001101011) && ({row_reg, col_reg}<20'b10001101010100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10001101010100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10001101010100011111) && ({row_reg, col_reg}<20'b10001101010101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10001101010101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10001101010101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10001101010101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10001101010101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10001101010101010000) && ({row_reg, col_reg}<20'b10001101011000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10001101011000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10001101011000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10001101011000111000) && ({row_reg, col_reg}<20'b10001101011000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10001101011000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10001101011000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10001101011000111100) && ({row_reg, col_reg}<20'b10001101011000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10001101011000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10001101011000111111) && ({row_reg, col_reg}<20'b10001101011001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10001101011001100110) && ({row_reg, col_reg}<20'b10001101011001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10001101011001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10001101011001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10001101011001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10001101011001101011) && ({row_reg, col_reg}<20'b10001101100100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10001101100100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10001101100100011111) && ({row_reg, col_reg}<20'b10001101100101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10001101100101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10001101100101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10001101100101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10001101100101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10001101100101010000) && ({row_reg, col_reg}<20'b10001101101000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10001101101000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10001101101000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10001101101000111000) && ({row_reg, col_reg}<20'b10001101101000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10001101101000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10001101101000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10001101101000111100) && ({row_reg, col_reg}<20'b10001101101000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10001101101000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10001101101000111111) && ({row_reg, col_reg}<20'b10001101101001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10001101101001100110) && ({row_reg, col_reg}<20'b10001101101001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10001101101001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10001101101001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10001101101001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10001101101001101011) && ({row_reg, col_reg}<20'b10001101110100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10001101110100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10001101110100011111) && ({row_reg, col_reg}<20'b10001101110101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10001101110101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10001101110101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10001101110101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10001101110101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10001101110101010000) && ({row_reg, col_reg}<20'b10001101111000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10001101111000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10001101111000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10001101111000111000) && ({row_reg, col_reg}<20'b10001101111000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10001101111000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10001101111000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10001101111000111100) && ({row_reg, col_reg}<20'b10001101111000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10001101111000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10001101111000111111) && ({row_reg, col_reg}<20'b10001101111001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10001101111001100110) && ({row_reg, col_reg}<20'b10001101111001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10001101111001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10001101111001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10001101111001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10001101111001101011) && ({row_reg, col_reg}<20'b10001110000100011001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=20'b10001110000100011001) && ({row_reg, col_reg}<20'b10001110000100011011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=20'b10001110000100011011) && ({row_reg, col_reg}<20'b10001110000100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10001110000100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10001110000100011111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10001110000100100000) && ({row_reg, col_reg}<20'b10001110000101001010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10001110000101001010) && ({row_reg, col_reg}<20'b10001110000101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10001110000101001100) && ({row_reg, col_reg}<20'b10001110000101001110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10001110000101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10001110000101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10001110000101010000) && ({row_reg, col_reg}<20'b10001110001000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10001110001000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10001110001000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==20'b10001110001000111000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10001110001000111001) && ({row_reg, col_reg}<20'b10001110001000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10001110001000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10001110001000111111) && ({row_reg, col_reg}<20'b10001110001001100001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10001110001001100001) && ({row_reg, col_reg}<20'b10001110001001100101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10001110001001100101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10001110001001100110) && ({row_reg, col_reg}<20'b10001110001001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10001110001001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10001110001001101001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=20'b10001110001001101010) && ({row_reg, col_reg}<20'b10001110001001101110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10001110001001101110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=20'b10001110001001101111) && ({row_reg, col_reg}<20'b10001110001101110000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10001110001101110000)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10001110001101110001) && ({row_reg, col_reg}<20'b10001110010100011100)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10001110010100011100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==20'b10001110010100011101)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10001110010100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10001110010100011111) && ({row_reg, col_reg}<20'b10001110010101001000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10001110010101001000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10001110010101001001) && ({row_reg, col_reg}<20'b10001110010101001110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10001110010101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10001110010101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10001110010101010000) && ({row_reg, col_reg}<20'b10001110011000110000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10001110011000110000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=20'b10001110011000110001) && ({row_reg, col_reg}<20'b10001110011000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10001110011000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10001110011000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10001110011000111000) && ({row_reg, col_reg}<20'b10001110011000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10001110011000111010) && ({row_reg, col_reg}<20'b10001110011000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10001110011000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10001110011000111111) && ({row_reg, col_reg}<20'b10001110011001100001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10001110011001100001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10001110011001100010) && ({row_reg, col_reg}<20'b10001110011001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10001110011001100110) && ({row_reg, col_reg}<20'b10001110011001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10001110011001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10001110011001101001) && ({row_reg, col_reg}<20'b10001110011001101100)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10001110011001101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=20'b10001110011001101101) && ({row_reg, col_reg}<20'b10001110011101101111)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10001110011101101111)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10001110011101110000) && ({row_reg, col_reg}<20'b10001110100100011100)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10001110100100011100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==20'b10001110100100011101)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10001110100100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10001110100100011111) && ({row_reg, col_reg}<20'b10001110100101001000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10001110100101001000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10001110100101001001) && ({row_reg, col_reg}<20'b10001110100101001011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10001110100101001011) && ({row_reg, col_reg}<20'b10001110100101001101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10001110100101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10001110100101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10001110100101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10001110100101010000) && ({row_reg, col_reg}<20'b10001110101000110000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10001110101000110000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=20'b10001110101000110001) && ({row_reg, col_reg}<20'b10001110101000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10001110101000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10001110101000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10001110101000111000) && ({row_reg, col_reg}<20'b10001110101000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10001110101000111010) && ({row_reg, col_reg}<20'b10001110101000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10001110101000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10001110101000111111) && ({row_reg, col_reg}<20'b10001110101001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10001110101001100110) && ({row_reg, col_reg}<20'b10001110101001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10001110101001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10001110101001101001) && ({row_reg, col_reg}<20'b10001110101001101100)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10001110101001101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=20'b10001110101001101101) && ({row_reg, col_reg}<20'b10001110101101101000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=20'b10001110101101101000) && ({row_reg, col_reg}<20'b10001110101101101011)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10001110101101101011) && ({row_reg, col_reg}<20'b10001110110000010000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=20'b10001110110000010000) && ({row_reg, col_reg}<20'b10001110110000010010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=20'b10001110110000010010) && ({row_reg, col_reg}<20'b10001110110100011000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=20'b10001110110100011000) && ({row_reg, col_reg}<20'b10001110110100011010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=20'b10001110110100011010) && ({row_reg, col_reg}<20'b10001110110100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10001110110100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10001110110100011111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10001110110100100000) && ({row_reg, col_reg}<20'b10001110110101001000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10001110110101001000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10001110110101001001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10001110110101001010) && ({row_reg, col_reg}<20'b10001110110101001101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10001110110101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10001110110101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10001110110101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10001110110101010000) && ({row_reg, col_reg}<20'b10001110110101010010)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10001110110101010010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=20'b10001110110101010011) && ({row_reg, col_reg}<20'b10001110111000110010)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10001110111000110010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=20'b10001110111000110011) && ({row_reg, col_reg}<20'b10001110111000110111)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10001110111000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10001110111000111000) && ({row_reg, col_reg}<20'b10001110111000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10001110111000111010) && ({row_reg, col_reg}<20'b10001110111000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10001110111000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10001110111000111111) && ({row_reg, col_reg}<20'b10001110111001100001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10001110111001100001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10001110111001100010) && ({row_reg, col_reg}<20'b10001110111001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10001110111001100110) && ({row_reg, col_reg}<20'b10001110111001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10001110111001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10001110111001101001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=20'b10001110111001101010) && ({row_reg, col_reg}<20'b10001110111001101100)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10001110111001101100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=20'b10001110111001101101) && ({row_reg, col_reg}<20'b10001110111001101111)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10001110111001101111)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10001110111001110000) && ({row_reg, col_reg}<20'b10001111000000010111)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10001111000000010111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=20'b10001111000000011000) && ({row_reg, col_reg}<20'b10001111000100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10001111000100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10001111000100011111) && ({row_reg, col_reg}<20'b10001111000101001000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10001111000101001000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10001111000101001001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10001111000101001010) && ({row_reg, col_reg}<20'b10001111000101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10001111000101001100) && ({row_reg, col_reg}<20'b10001111000101001110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10001111000101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10001111000101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10001111000101010000) && ({row_reg, col_reg}<20'b10001111001000110010)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10001111001000110010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=20'b10001111001000110011) && ({row_reg, col_reg}<20'b10001111001000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10001111001000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10001111001000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10001111001000111000) && ({row_reg, col_reg}<20'b10001111001000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10001111001000111010) && ({row_reg, col_reg}<20'b10001111001000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10001111001000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10001111001000111111) && ({row_reg, col_reg}<20'b10001111001001100000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10001111001001100000) && ({row_reg, col_reg}<20'b10001111001001100010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10001111001001100010) && ({row_reg, col_reg}<20'b10001111001001100100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10001111001001100100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10001111001001100101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10001111001001100110) && ({row_reg, col_reg}<20'b10001111001001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10001111001001101000)) color_data = 12'b101110111011;

		if(({row_reg, col_reg}>=20'b10001111001001101001) && ({row_reg, col_reg}<20'b10001111010000001110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=20'b10001111010000001110) && ({row_reg, col_reg}<20'b10001111010000010000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=20'b10001111010000010000) && ({row_reg, col_reg}<20'b10001111010000011000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=20'b10001111010000011000) && ({row_reg, col_reg}<20'b10001111010000011010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=20'b10001111010000011010) && ({row_reg, col_reg}<20'b10001111010100011100)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10001111010100011100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==20'b10001111010100011101)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10001111010100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10001111010100011111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10001111010100100000) && ({row_reg, col_reg}<20'b10001111010101001000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10001111010101001000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10001111010101001001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10001111010101001010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10001111010101001011) && ({row_reg, col_reg}<20'b10001111010101001110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10001111010101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10001111010101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10001111010101010000) && ({row_reg, col_reg}<20'b10001111010101010100)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10001111010101010100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=20'b10001111010101010101) && ({row_reg, col_reg}<20'b10001111011000110100)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=20'b10001111011000110100) && ({row_reg, col_reg}<20'b10001111011000110110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==20'b10001111011000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10001111011000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10001111011000111000) && ({row_reg, col_reg}<20'b10001111011000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10001111011000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10001111011000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10001111011000111100) && ({row_reg, col_reg}<20'b10001111011000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10001111011000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10001111011000111111) && ({row_reg, col_reg}<20'b10001111011001100000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10001111011001100000) && ({row_reg, col_reg}<20'b10001111011001100010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10001111011001100010) && ({row_reg, col_reg}<20'b10001111011001100100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10001111011001100100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10001111011001100101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10001111011001100110) && ({row_reg, col_reg}<20'b10001111011001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10001111011001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10001111011001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10001111011001101010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=20'b10001111011001101011) && ({row_reg, col_reg}<20'b10001111011001101101)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10001111011001101101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=20'b10001111011001101110) && ({row_reg, col_reg}<20'b10001111011101101111)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10001111011101101111)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10001111011101110000) && ({row_reg, col_reg}<20'b10001111100000010101)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=20'b10001111100000010101) && ({row_reg, col_reg}<20'b10001111100000011000)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=20'b10001111100000011000) && ({row_reg, col_reg}<20'b10001111100100011110)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==20'b10001111100100011110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=20'b10001111100100011111) && ({row_reg, col_reg}<20'b10001111100101001010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10001111100101001010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10001111100101001011) && ({row_reg, col_reg}<20'b10001111100101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10001111100101001101) && ({row_reg, col_reg}<20'b10001111100101001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10001111100101001111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==20'b10001111100101010000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10001111100101010001) && ({row_reg, col_reg}<20'b10001111101000110110)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==20'b10001111101000110110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10001111101000110111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==20'b10001111101000111000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10001111101000111001) && ({row_reg, col_reg}<20'b10001111101000111011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10001111101000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10001111101000111100) && ({row_reg, col_reg}<20'b10001111101001100100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10001111101001100100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10001111101001100101) && ({row_reg, col_reg}<20'b10001111101001100111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10001111101001100111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10001111101001101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10001111101001101001) && ({row_reg, col_reg}<20'b10001111101101101010)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=20'b10001111101101101010) && ({row_reg, col_reg}<20'b10001111101101101101)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=20'b10001111101101101101) && ({row_reg, col_reg}<20'b10001111101101101111)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10001111101101101111)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10001111101101110000) && ({row_reg, col_reg}<20'b10001111110000010001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=20'b10001111110000010001) && ({row_reg, col_reg}<20'b10001111110000010100)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10001111110000010100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==20'b10001111110000010101)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10001111110000010110) && ({row_reg, col_reg}<20'b10001111110000011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10001111110000011000) && ({row_reg, col_reg}<20'b10001111110100011110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=20'b10001111110100011110) && ({row_reg, col_reg}<20'b10001111110100100000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10001111110100100000) && ({row_reg, col_reg}<20'b10001111110101001010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10001111110101001010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10001111110101001011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10001111110101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10001111110101001101) && ({row_reg, col_reg}<20'b10001111110101001111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10001111110101001111) && ({row_reg, col_reg}<20'b10001111110101010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10001111110101010001) && ({row_reg, col_reg}<20'b10001111111000110101)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==20'b10001111111000110101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10001111111000110110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=20'b10001111111000110111) && ({row_reg, col_reg}<20'b10001111111000111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10001111111000111001) && ({row_reg, col_reg}<20'b10001111111000111011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10001111111000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10001111111000111100) && ({row_reg, col_reg}<20'b10001111111001100100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10001111111001100100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10001111111001100101) && ({row_reg, col_reg}<20'b10001111111001100111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10001111111001100111) && ({row_reg, col_reg}<20'b10001111111001101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10001111111001101001) && ({row_reg, col_reg}<20'b10001111111101101010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==20'b10001111111101101010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10001111111101101011) && ({row_reg, col_reg}<20'b10001111111101101101)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10001111111101101101)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=20'b10001111111101101110) && ({row_reg, col_reg}<20'b10001111111101110000)) color_data = 12'b110111011101;

		if(({row_reg, col_reg}>=20'b10001111111101110000) && ({row_reg, col_reg}<20'b10010000000000001001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=20'b10010000000000001001) && ({row_reg, col_reg}<20'b10010000000000001011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=20'b10010000000000001011) && ({row_reg, col_reg}<20'b10010000000000001110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10010000000000001110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10010000000000001111)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10010000000000010000) && ({row_reg, col_reg}<20'b10010000000000010010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10010000000000010010) && ({row_reg, col_reg}<20'b10010000000000010100)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=20'b10010000000000010100) && ({row_reg, col_reg}<20'b10010000000100100000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10010000000100100000) && ({row_reg, col_reg}<20'b10010000000101010000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10010000000101010000) && ({row_reg, col_reg}<20'b10010000001000111000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10010000001000111000) && ({row_reg, col_reg}<20'b10010000001001101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10010000001001101000) && ({row_reg, col_reg}<20'b10010000001101101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10010000001101101110) && ({row_reg, col_reg}<20'b10010000001101110000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==20'b10010000001101110000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==20'b10010000001101110001)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10010000001101110010)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=20'b10010000001101110011) && ({row_reg, col_reg}<20'b10010000001101111010)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10010000001101111010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=20'b10010000001101111011) && ({row_reg, col_reg}<20'b10010000001101111101)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=20'b10010000001101111101) && ({row_reg, col_reg}<20'b10010000001101111111)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10010000001101111111) && ({row_reg, col_reg}<20'b10010000010000001010)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10010000010000001010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==20'b10010000010000001011)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10010000010000001100)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10010000010000001101)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==20'b10010000010000001110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==20'b10010000010000001111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=20'b10010000010000010000) && ({row_reg, col_reg}<20'b10010000010000010011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10010000010000010011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10010000010000010100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10010000010000010101) && ({row_reg, col_reg}<20'b10010000011101101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10010000011101101101) && ({row_reg, col_reg}<20'b10010000011101110001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10010000011101110001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==20'b10010000011101110010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==20'b10010000011101110011)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==20'b10010000011101110100)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=20'b10010000011101110101) && ({row_reg, col_reg}<20'b10010000011101110111)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10010000011101110111)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10010000011101111000) && ({row_reg, col_reg}<20'b10010000100000000011)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10010000100000000011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=20'b10010000100000000100) && ({row_reg, col_reg}<20'b10010000100000001000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10010000100000001000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=20'b10010000100000001001) && ({row_reg, col_reg}<20'b10010000100000001011)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10010000100000001011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10010000100000001100)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10010000100000001101)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=20'b10010000100000001110) && ({row_reg, col_reg}<20'b10010000100000010000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10010000100000010000) && ({row_reg, col_reg}<20'b10010000100000010111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10010000100000010111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10010000100000011000) && ({row_reg, col_reg}<20'b10010000101101110010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10010000101101110010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10010000101101110011)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==20'b10010000101101110100)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10010000101101110101)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=20'b10010000101101110110) && ({row_reg, col_reg}<20'b10010000101101111000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10010000101101111000)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10010000101101111001) && ({row_reg, col_reg}<20'b10010000110000001000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10010000110000001000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==20'b10010000110000001001)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10010000110000001010)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==20'b10010000110000001011)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10010000110000001100) && ({row_reg, col_reg}<20'b10010000110000001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10010000110000001110) && ({row_reg, col_reg}<20'b10010000110000010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10010000110000010001) && ({row_reg, col_reg}<20'b10010000110000010101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10010000110000010101) && ({row_reg, col_reg}<20'b10010000111101101110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10010000111101101110) && ({row_reg, col_reg}<20'b10010000111101110001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10010000111101110001) && ({row_reg, col_reg}<20'b10010000111101110011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10010000111101110011) && ({row_reg, col_reg}<20'b10010000111101110101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10010000111101110101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==20'b10010000111101110110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10010000111101110111)) color_data = 12'b110111011101;

		if(({row_reg, col_reg}>=20'b10010000111101111000) && ({row_reg, col_reg}<20'b10010001000000000101)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10010001000000000101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=20'b10010001000000000110) && ({row_reg, col_reg}<20'b10010001000000001000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10010001000000001000)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10010001000000001001)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10010001000000001010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==20'b10010001000000001011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10010001000000001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10010001000000001101) && ({row_reg, col_reg}<20'b10010001000000001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10010001000000001111) && ({row_reg, col_reg}<20'b10010001001101110010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10010001001101110010) && ({row_reg, col_reg}<20'b10010001001101110100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10010001001101110100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10010001001101110101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10010001001101110110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==20'b10010001001101110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==20'b10010001001101111000)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=20'b10010001001101111001) && ({row_reg, col_reg}<20'b10010001010000000001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10010001010000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=20'b10010001010000000010) && ({row_reg, col_reg}<20'b10010001010000000101)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10010001010000000101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==20'b10010001010000000110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10010001010000000111)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==20'b10010001010000001000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==20'b10010001010000001001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10010001010000001010) && ({row_reg, col_reg}<20'b10010001010000001111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10010001010000001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10010001010000010000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10010001010000010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10010001010000010010) && ({row_reg, col_reg}<20'b10010001010000010100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10010001010000010100) && ({row_reg, col_reg}<20'b10010001010000011000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10010001010000011000) && ({row_reg, col_reg}<20'b10010001011101101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10010001011101101000) && ({row_reg, col_reg}<20'b10010001011101101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10010001011101101110) && ({row_reg, col_reg}<20'b10010001011101110000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10010001011101110000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10010001011101110001) && ({row_reg, col_reg}<20'b10010001011101110100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10010001011101110100) && ({row_reg, col_reg}<20'b10010001011101111000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10010001011101111000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==20'b10010001011101111001)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=20'b10010001011101111010) && ({row_reg, col_reg}<20'b10010001100000000110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10010001100000000110)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==20'b10010001100000000111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==20'b10010001100000001000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10010001100000001001) && ({row_reg, col_reg}<20'b10010001100000001011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10010001100000001011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10010001100000001100) && ({row_reg, col_reg}<20'b10010001100000001111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10010001100000001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10010001100000010000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10010001100000010001) && ({row_reg, col_reg}<20'b10010001100000010011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10010001100000010011) && ({row_reg, col_reg}<20'b10010001101101110001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10010001101101110001) && ({row_reg, col_reg}<20'b10010001101101110100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10010001101101110100) && ({row_reg, col_reg}<20'b10010001101101110111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10010001101101110111) && ({row_reg, col_reg}<20'b10010001101101111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10010001101101111001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==20'b10010001101101111010)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=20'b10010001101101111011) && ({row_reg, col_reg}<20'b10010001110000000101)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10010001110000000101)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10010001110000000110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==20'b10010001110000000111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10010001110000001000) && ({row_reg, col_reg}<20'b10010001110000001010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10010001110000001010) && ({row_reg, col_reg}<20'b10010001110000001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10010001110000001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10010001110000001101) && ({row_reg, col_reg}<20'b10010001110000001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10010001110000001111) && ({row_reg, col_reg}<20'b10010001110000010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10010001110000010001) && ({row_reg, col_reg}<20'b10010001110000010100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10010001110000010100) && ({row_reg, col_reg}<20'b10010001110000010110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10010001110000010110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10010001110000010111) && ({row_reg, col_reg}<20'b10010001111101101001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10010001111101101001) && ({row_reg, col_reg}<20'b10010001111101101101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10010001111101101101) && ({row_reg, col_reg}<20'b10010001111101110100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10010001111101110100) && ({row_reg, col_reg}<20'b10010001111101110110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10010001111101110110) && ({row_reg, col_reg}<20'b10010001111101111000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10010001111101111000) && ({row_reg, col_reg}<20'b10010001111101111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10010001111101111010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==20'b10010001111101111011)) color_data = 12'b110111011101;

		if(({row_reg, col_reg}>=20'b10010001111101111100) && ({row_reg, col_reg}<20'b10010010000000000100)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10010010000000000100)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10010010000000000101)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10010010000000000110) && ({row_reg, col_reg}<20'b10010010000000001000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10010010000000001000) && ({row_reg, col_reg}<20'b10010010001101111000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10010010001101111000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10010010001101111001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10010010001101111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10010010001101111011)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10010010001101111100)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10010010001101111101)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10010010001101111110) && ({row_reg, col_reg}<20'b10010010010000000010)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10010010010000000010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==20'b10010010010000000011)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10010010010000000100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==20'b10010010010000000101)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=20'b10010010010000000110) && ({row_reg, col_reg}<20'b10010010010000001000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10010010010000001000) && ({row_reg, col_reg}<20'b10010010011101111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10010010011101111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10010010011101111011)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==20'b10010010011101111100)) color_data = 12'b101110111011;

		if(({row_reg, col_reg}>=20'b10010010011101111101) && ({row_reg, col_reg}<20'b10010010100000000011)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10010010100000000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10010010100000000100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10010010100000000101) && ({row_reg, col_reg}<20'b10010010100000000111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10010010100000000111) && ({row_reg, col_reg}<20'b10010010101101111001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10010010101101111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10010010101101111010) && ({row_reg, col_reg}<20'b10010010101101111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10010010101101111100)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==20'b10010010101101111101)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=20'b10010010101101111110) && ({row_reg, col_reg}<20'b10010010110000000010)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10010010110000000010)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10010010110000000011)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10010010110000000100)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=20'b10010010110000000101) && ({row_reg, col_reg}<20'b10010010110000000111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10010010110000000111) && ({row_reg, col_reg}<20'b10010010111101111001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10010010111101111001) && ({row_reg, col_reg}<20'b10010010111101111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10010010111101111011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10010010111101111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10010010111101111101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==20'b10010010111101111110)) color_data = 12'b110111011101;

		if(({row_reg, col_reg}>=20'b10010010111101111111) && ({row_reg, col_reg}<20'b10010011000000000010)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10010011000000000010)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10010011000000000011)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==20'b10010011000000000100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10010011000000000101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10010011000000000110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10010011000000000111) && ({row_reg, col_reg}<20'b10010011001101111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10010011001101111010) && ({row_reg, col_reg}<20'b10010011001101111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10010011001101111110)) color_data = 12'b101110111011;

		if(({row_reg, col_reg}>=20'b10010011001101111111) && ({row_reg, col_reg}<20'b10010011010000000001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10010011010000000001)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10010011010000000010)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10010011010000000011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10010011010000000100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10010011010000000101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10010011010000000110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10010011010000000111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10010011010000001000) && ({row_reg, col_reg}<20'b10010011011101111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10010011011101111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10010011011101111011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10010011011101111100) && ({row_reg, col_reg}<20'b10010011011101111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10010011011101111110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==20'b10010011011101111111)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=20'b10010011011110000000) && ({row_reg, col_reg}<20'b10010011100000000001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10010011100000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==20'b10010011100000000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=20'b10010011100000000011) && ({row_reg, col_reg}<20'b10010011100000000110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10010011100000000110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10010011100000000111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10010011100000001000) && ({row_reg, col_reg}<20'b10010011101101111000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10010011101101111000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10010011101101111001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10010011101101111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10010011101101111011) && ({row_reg, col_reg}<20'b10010011101101111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10010011101101111101) && ({row_reg, col_reg}<20'b10010011101101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10010011101101111111)) color_data = 12'b101110111011;

		if(({row_reg, col_reg}>=20'b10010011101110000000) && ({row_reg, col_reg}<20'b10010011110000000001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10010011110000000001)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10010011110000000010) && ({row_reg, col_reg}<20'b10010011110000000100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10010011110000000100) && ({row_reg, col_reg}<20'b10010011110000000110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10010011110000000110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10010011110000000111) && ({row_reg, col_reg}<20'b10010011111101111000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10010011111101111000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10010011111101111001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10010011111101111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10010011111101111011) && ({row_reg, col_reg}<20'b10010011111101111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10010011111101111101) && ({row_reg, col_reg}<20'b10010011111101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10010011111101111111)) color_data = 12'b101110111011;

		if(({row_reg, col_reg}>=20'b10010011111110000000) && ({row_reg, col_reg}<20'b10010100000000000001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10010100000000000001)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10010100000000000010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10010100000000000011) && ({row_reg, col_reg}<20'b10010100000000000101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10010100000000000101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10010100000000000110) && ({row_reg, col_reg}<20'b10010100001101111000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10010100001101111000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10010100001101111001) && ({row_reg, col_reg}<20'b10010100001101111011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10010100001101111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10010100001101111100) && ({row_reg, col_reg}<20'b10010100001101111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10010100001101111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10010100001101111111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==20'b10010100001110000000)) color_data = 12'b110111011101;

		if(({row_reg, col_reg}>=20'b10010100001110000001) && ({row_reg, col_reg}<20'b10010100010000000000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10010100010000000000)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10010100010000000001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==20'b10010100010000000010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10010100010000000011) && ({row_reg, col_reg}<20'b10010100011101111000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10010100011101111000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10010100011101111001) && ({row_reg, col_reg}<20'b10010100011101111011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10010100011101111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10010100011101111100) && ({row_reg, col_reg}<20'b10010100011101111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10010100011101111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10010100011101111111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==20'b10010100011110000000)) color_data = 12'b110111011101;

		if(({row_reg, col_reg}>=20'b10010100011110000001) && ({row_reg, col_reg}<20'b10010100100000000000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10010100100000000000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==20'b10010100100000000001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10010100100000000010) && ({row_reg, col_reg}<20'b10010100100000000100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10010100100000000100) && ({row_reg, col_reg}<20'b10010100100000000111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10010100100000000111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10010100100000001000) && ({row_reg, col_reg}<20'b10010100101101111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10010100101101111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10010100101101111011) && ({row_reg, col_reg}<20'b10010100101101111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10010100101101111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10010100101101111111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==20'b10010100101110000000)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=20'b10010100101110000001) && ({row_reg, col_reg}<20'b10010100110000000000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10010100110000000000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10010100110000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==20'b10010100110000000010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10010100110000000011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10010100110000000100) && ({row_reg, col_reg}<20'b10010100111101111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10010100111101111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10010100111101111011) && ({row_reg, col_reg}<20'b10010100111101111111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10010100111101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10010100111110000000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10010100111110000001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10010100111110000010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}==20'b10010100111110000011)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10010101000000000000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==20'b10010101000000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==20'b10010101000000000010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10010101000000000011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10010101000000000100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10010101000000000101) && ({row_reg, col_reg}<20'b10010101000000000111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10010101000000000111) && ({row_reg, col_reg}<20'b10010101001101111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10010101001101111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10010101001101111011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10010101001101111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10010101001101111101) && ({row_reg, col_reg}<20'b10010101001101111111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10010101001101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10010101001110000000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==20'b10010101001110000001)) color_data = 12'b110111011101;

		if(({row_reg, col_reg}>=20'b10010101001110000010) && ({row_reg, col_reg}<20'b10010101010000000000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==20'b10010101010000000000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==20'b10010101010000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==20'b10010101010000000010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10010101010000000011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10010101010000000100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10010101010000000101) && ({row_reg, col_reg}<20'b10010101010000000111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10010101010000000111) && ({row_reg, col_reg}<20'b10010101011101111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10010101011101111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10010101011101111011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10010101011101111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10010101011101111101) && ({row_reg, col_reg}<20'b10010101011101111111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10010101011101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10010101011110000000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==20'b10010101011110000001)) color_data = 12'b110111011101;

		if(({row_reg, col_reg}>=20'b10010101011110000010) && ({row_reg, col_reg}<20'b10010101100000000000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10010101100000000000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==20'b10010101100000000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10010101100000000010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10010101100000000011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10010101100000000100) && ({row_reg, col_reg}<20'b10010101100000000110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10010101100000000110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10010101100000000111) && ({row_reg, col_reg}<20'b10010101101101111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10010101101101111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10010101101101111011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10010101101101111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10010101101101111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10010101101101111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10010101101101111111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10010101101110000000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==20'b10010101101110000001)) color_data = 12'b110111011101;

		if(({row_reg, col_reg}>=20'b10010101101110000010) && ({row_reg, col_reg}<20'b10010101110000000000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=20'b10010101110000000000) && ({row_reg, col_reg}<20'b10010101110000000010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10010101110000000010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10010101110000000011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10010101110000000100) && ({row_reg, col_reg}<20'b10010101110000000110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10010101110000000110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10010101110000000111) && ({row_reg, col_reg}<20'b10010101111101111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10010101111101111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10010101111101111011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10010101111101111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10010101111101111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10010101111101111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10010101111101111111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10010101111110000000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==20'b10010101111110000001)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10010101111110000010)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}==20'b10010101111110000011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=20'b10010110000000000000) && ({row_reg, col_reg}<20'b10010110000000000010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10010110000000000010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10010110000000000011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10010110000000000100) && ({row_reg, col_reg}<20'b10010110000000000110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10010110000000000110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10010110000000000111) && ({row_reg, col_reg}<20'b10010110001101111001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10010110001101111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10010110001101111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10010110001101111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10010110001101111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10010110001101111101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10010110001101111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10010110001101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10010110001110000000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==20'b10010110001110000001)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10010110001110000010)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}==20'b10010110001110000011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==20'b10010110010000000000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==20'b10010110010000000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10010110010000000010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10010110010000000011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10010110010000000100) && ({row_reg, col_reg}<20'b10010110010000000110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10010110010000000110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10010110010000000111) && ({row_reg, col_reg}<20'b10010110011101111001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10010110011101111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10010110011101111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10010110011101111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10010110011101111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10010110011101111101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10010110011101111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10010110011101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10010110011110000000)) color_data = 12'b101010101010;

		if(({row_reg, col_reg}>=20'b10010110011110000001) && ({row_reg, col_reg}<20'b10010110100000000000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10010110100000000000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==20'b10010110100000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==20'b10010110100000000010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10010110100000000011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10010110100000000100) && ({row_reg, col_reg}<20'b10010110101101111001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10010110101101111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10010110101101111010) && ({row_reg, col_reg}<20'b10010110101101111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10010110101101111101) && ({row_reg, col_reg}<20'b10010110101110000000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10010110101110000000)) color_data = 12'b101110111011;

		if(({row_reg, col_reg}>=20'b10010110101110000001) && ({row_reg, col_reg}<20'b10010110110000000000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10010110110000000000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10010110110000000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==20'b10010110110000000010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10010110110000000011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10010110110000000100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10010110110000000101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10010110110000000110) && ({row_reg, col_reg}<20'b10010110111101111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10010110111101111101) && ({row_reg, col_reg}<20'b10010110111101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10010110111101111111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==20'b10010110111110000000)) color_data = 12'b101110111011;

		if(({row_reg, col_reg}>=20'b10010110111110000001) && ({row_reg, col_reg}<20'b10010111000000000000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10010111000000000000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==20'b10010111000000000001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10010111000000000010) && ({row_reg, col_reg}<20'b10010111000000000101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10010111000000000101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10010111000000000110) && ({row_reg, col_reg}<20'b10010111001101111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10010111001101111010) && ({row_reg, col_reg}<20'b10010111001101111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10010111001101111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10010111001101111101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10010111001101111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10010111001101111111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==20'b10010111001110000000)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=20'b10010111001110000001) && ({row_reg, col_reg}<20'b10010111010000000000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10010111010000000000)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10010111010000000001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==20'b10010111010000000010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10010111010000000011) && ({row_reg, col_reg}<20'b10010111010000000101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10010111010000000101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10010111010000000110) && ({row_reg, col_reg}<20'b10010111011101111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10010111011101111010) && ({row_reg, col_reg}<20'b10010111011101111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10010111011101111100) && ({row_reg, col_reg}<20'b10010111011101111111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10010111011101111111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==20'b10010111011110000000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=20'b10010111011110000001) && ({row_reg, col_reg}<20'b10010111011110000011)) color_data = 12'b111011101110;

		if(({row_reg, col_reg}==20'b10010111011110000011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==20'b10010111100000000000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10010111100000000001)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10010111100000000010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10010111100000000011) && ({row_reg, col_reg}<20'b10010111100000000101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10010111100000000101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10010111100000000110) && ({row_reg, col_reg}<20'b10010111101101111000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10010111101101111000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10010111101101111001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10010111101101111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10010111101101111011) && ({row_reg, col_reg}<20'b10010111101101111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10010111101101111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10010111101101111111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==20'b10010111101110000000)) color_data = 12'b110111011101;

		if(({row_reg, col_reg}>=20'b10010111101110000001) && ({row_reg, col_reg}<20'b10010111110000000000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10010111110000000000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==20'b10010111110000000001)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10010111110000000010) && ({row_reg, col_reg}<20'b10010111110000000100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10010111110000000100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10010111110000000101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10010111110000000110) && ({row_reg, col_reg}<20'b10010111111101111000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10010111111101111000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10010111111101111001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10010111111101111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10010111111101111011) && ({row_reg, col_reg}<20'b10010111111101111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10010111111101111101) && ({row_reg, col_reg}<20'b10010111111101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10010111111101111111)) color_data = 12'b101110111011;

		if(({row_reg, col_reg}>=20'b10010111111110000000) && ({row_reg, col_reg}<20'b10011000000000000001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10011000000000000001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==20'b10011000000000000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==20'b10011000000000000011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10011000000000000100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10011000000000000101) && ({row_reg, col_reg}<20'b10011000000000000111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10011000000000000111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10011000000000001000) && ({row_reg, col_reg}<20'b10011000001101111001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10011000001101111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10011000001101111010) && ({row_reg, col_reg}<20'b10011000001101111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10011000001101111101) && ({row_reg, col_reg}<20'b10011000001101111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10011000001101111111)) color_data = 12'b101110111011;

		if(({row_reg, col_reg}>=20'b10011000001110000000) && ({row_reg, col_reg}<20'b10011000010000000001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10011000010000000001)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10011000010000000010)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10011000010000000011) && ({row_reg, col_reg}<20'b10011000010000000101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10011000010000000101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10011000010000000110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10011000010000000111) && ({row_reg, col_reg}<20'b10011000011101111000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10011000011101111000) && ({row_reg, col_reg}<20'b10011000011101111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10011000011101111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10011000011101111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10011000011101111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10011000011101111101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10011000011101111110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==20'b10011000011101111111)) color_data = 12'b110111011101;

		if(({row_reg, col_reg}>=20'b10011000011110000000) && ({row_reg, col_reg}<20'b10011000100000000010)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10011000100000000010)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==20'b10011000100000000011)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==20'b10011000100000000100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10011000100000000101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10011000100000000110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10011000100000000111) && ({row_reg, col_reg}<20'b10011000101101111000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10011000101101111000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10011000101101111001) && ({row_reg, col_reg}<20'b10011000101101111011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10011000101101111011) && ({row_reg, col_reg}<20'b10011000101101111101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10011000101101111101)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==20'b10011000101101111110)) color_data = 12'b110111011101;

		if(({row_reg, col_reg}>=20'b10011000101101111111) && ({row_reg, col_reg}<20'b10011000110000000001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10011000110000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==20'b10011000110000000010)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10011000110000000011)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10011000110000000100)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==20'b10011000110000000101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10011000110000000110) && ({row_reg, col_reg}<20'b10011000111101111000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10011000111101111000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10011000111101111001) && ({row_reg, col_reg}<20'b10011000111101111011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10011000111101111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10011000111101111100)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==20'b10011000111101111101)) color_data = 12'b101110111011;

		if(({row_reg, col_reg}>=20'b10011000111101111110) && ({row_reg, col_reg}<20'b10011001000000000011)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10011001000000000011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10011001000000000100)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10011001000000000101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10011001000000000110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10011001000000000111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10011001000000001000) && ({row_reg, col_reg}<20'b10011001001101111000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10011001001101111000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10011001001101111001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10011001001101111010) && ({row_reg, col_reg}<20'b10011001001101111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10011001001101111100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==20'b10011001001101111101)) color_data = 12'b110111011101;

		if(({row_reg, col_reg}>=20'b10011001001101111110) && ({row_reg, col_reg}<20'b10011001010000000100)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10011001010000000100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==20'b10011001010000000101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==20'b10011001010000000110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10011001010000000111) && ({row_reg, col_reg}<20'b10011001011101111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10011001011101111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10011001011101111011)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==20'b10011001011101111100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=20'b10011001011101111101) && ({row_reg, col_reg}<20'b10011001100000000001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10011001100000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==20'b10011001100000000010)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10011001100000000011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==20'b10011001100000000100)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10011001100000000101)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==20'b10011001100000000110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==20'b10011001100000000111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10011001100000001000) && ({row_reg, col_reg}<20'b10011001101101111001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10011001101101111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10011001101101111010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==20'b10011001101101111011)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10011001101101111100)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10011001101101111101)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10011001101101111110) && ({row_reg, col_reg}<20'b10011001110000000001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10011001110000000001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=20'b10011001110000000010) && ({row_reg, col_reg}<20'b10011001110000000100)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10011001110000000100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==20'b10011001110000000101)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10011001110000000110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10011001110000000111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=20'b10011001110000001000) && ({row_reg, col_reg}<20'b10011001111101111001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10011001111101111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10011001111101111010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==20'b10011001111101111011)) color_data = 12'b110111011101;

		if(({row_reg, col_reg}>=20'b10011001111101111100) && ({row_reg, col_reg}<20'b10011010000000000110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10011010000000000110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10011010000000000111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10011010000000001000) && ({row_reg, col_reg}<20'b10011010000000001010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10011010000000001010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10011010000000001011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10011010000000001100) && ({row_reg, col_reg}<20'b10011010000000001111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10011010000000001111) && ({row_reg, col_reg}<20'b10011010000000010010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10011010000000010010) && ({row_reg, col_reg}<20'b10011010000100011011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10011010000100011011) && ({row_reg, col_reg}<20'b10011010000100011101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10011010000100011101) && ({row_reg, col_reg}<20'b10011010000101001000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10011010000101001000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10011010000101001001) && ({row_reg, col_reg}<20'b10011010000101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10011010000101001100) && ({row_reg, col_reg}<20'b10011010000101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10011010000101001110) && ({row_reg, col_reg}<20'b10011010001000110000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10011010001000110000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10011010001000110001) && ({row_reg, col_reg}<20'b10011010001001101001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10011010001001101001) && ({row_reg, col_reg}<20'b10011010001001101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10011010001001101100) && ({row_reg, col_reg}<20'b10011010001001101111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10011010001001101111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10011010001001110000) && ({row_reg, col_reg}<20'b10011010001101110001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10011010001101110001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10011010001101110010) && ({row_reg, col_reg}<20'b10011010001101110101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10011010001101110101) && ({row_reg, col_reg}<20'b10011010001101110111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10011010001101110111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10011010001101111000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10011010001101111001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==20'b10011010001101111010)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==20'b10011010001101111011)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10011010001101111100)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10011010001101111101) && ({row_reg, col_reg}<20'b10011010010000000101)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10011010010000000101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==20'b10011010010000000110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10011010010000000111)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==20'b10011010010000001000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==20'b10011010010000001001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==20'b10011010010000001010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10011010010000001011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10011010010000001100) && ({row_reg, col_reg}<20'b10011010010000001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10011010010000001111) && ({row_reg, col_reg}<20'b10011010010100011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10011010010100011000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10011010010100011001) && ({row_reg, col_reg}<20'b10011010010101001000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10011010010101001000) && ({row_reg, col_reg}<20'b10011010010101001010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10011010010101001010) && ({row_reg, col_reg}<20'b10011010011000110000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10011010011000110000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10011010011000110001) && ({row_reg, col_reg}<20'b10011010011000110011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10011010011000110011) && ({row_reg, col_reg}<20'b10011010011000111000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10011010011000111000) && ({row_reg, col_reg}<20'b10011010011101101011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10011010011101101011) && ({row_reg, col_reg}<20'b10011010011101110001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10011010011101110001) && ({row_reg, col_reg}<20'b10011010011101110011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10011010011101110011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10011010011101110100) && ({row_reg, col_reg}<20'b10011010011101110110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10011010011101110110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10011010011101110111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==20'b10011010011101111000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==20'b10011010011101111001)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=20'b10011010011101111010) && ({row_reg, col_reg}<20'b10011010100000000000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10011010100000000000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=20'b10011010100000000001) && ({row_reg, col_reg}<20'b10011010100000000101)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=20'b10011010100000000101) && ({row_reg, col_reg}<20'b10011010100000000111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==20'b10011010100000000111)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10011010100000001000)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10011010100000001001)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10011010100000001010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==20'b10011010100000001011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10011010100000001100) && ({row_reg, col_reg}<20'b10011010100000001110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10011010100000001110) && ({row_reg, col_reg}<20'b10011010100000010000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10011010100000010000) && ({row_reg, col_reg}<20'b10011010100000010100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10011010100000010100) && ({row_reg, col_reg}<20'b10011010100000011000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10011010100000011000) && ({row_reg, col_reg}<20'b10011010100100011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10011010100100011000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10011010100100011001) && ({row_reg, col_reg}<20'b10011010100100011101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10011010100100011101) && ({row_reg, col_reg}<20'b10011010100100100000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10011010100100100000) && ({row_reg, col_reg}<20'b10011010100101001000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10011010100101001000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10011010100101001001) && ({row_reg, col_reg}<20'b10011010101101101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10011010101101101000) && ({row_reg, col_reg}<20'b10011010101101101010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10011010101101101010) && ({row_reg, col_reg}<20'b10011010101101110000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10011010101101110000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10011010101101110001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10011010101101110010) && ({row_reg, col_reg}<20'b10011010101101110100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10011010101101110100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10011010101101110101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10011010101101110110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==20'b10011010101101110111)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==20'b10011010101101111000)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10011010101101111001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=20'b10011010101101111010) && ({row_reg, col_reg}<20'b10011010101101111100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=20'b10011010101101111100) && ({row_reg, col_reg}<20'b10011010101101111110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10011010101101111110)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10011010101101111111) && ({row_reg, col_reg}<20'b10011010110000001000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10011010110000001000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==20'b10011010110000001001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10011010110000001010)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==20'b10011010110000001011)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10011010110000001100)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==20'b10011010110000001101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10011010110000001110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10011010110000001111) && ({row_reg, col_reg}<20'b10011010110000010101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10011010110000010101) && ({row_reg, col_reg}<20'b10011010110000011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10011010110000011000) && ({row_reg, col_reg}<20'b10011010110000011010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10011010110000011010) && ({row_reg, col_reg}<20'b10011010110000011101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10011010110000011101) && ({row_reg, col_reg}<20'b10011010110000100000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10011010110000100000) && ({row_reg, col_reg}<20'b10011010110101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10011010110101001100) && ({row_reg, col_reg}<20'b10011010110101010000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10011010110101010000) && ({row_reg, col_reg}<20'b10011010111000110000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10011010111000110000) && ({row_reg, col_reg}<20'b10011010111000111000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10011010111000111000) && ({row_reg, col_reg}<20'b10011010111001101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10011010111001101000) && ({row_reg, col_reg}<20'b10011010111001101010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10011010111001101010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10011010111001101011) && ({row_reg, col_reg}<20'b10011010111001110000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10011010111001110000) && ({row_reg, col_reg}<20'b10011010111101101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10011010111101101100) && ({row_reg, col_reg}<20'b10011010111101110001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10011010111101110001) && ({row_reg, col_reg}<20'b10011010111101110011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10011010111101110011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10011010111101110100)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==20'b10011010111101110101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==20'b10011010111101110110)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=20'b10011010111101110111) && ({row_reg, col_reg}<20'b10011011000000000011)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10011011000000000011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=20'b10011011000000000100) && ({row_reg, col_reg}<20'b10011011000000001100)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10011011000000001100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==20'b10011011000000001101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==20'b10011011000000001110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==20'b10011011000000001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10011011000000010000) && ({row_reg, col_reg}<20'b10011011000000010110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10011011000000010110) && ({row_reg, col_reg}<20'b10011011000000011000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10011011000000011000) && ({row_reg, col_reg}<20'b10011011000100011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10011011000100011000) && ({row_reg, col_reg}<20'b10011011000100011101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10011011000100011101) && ({row_reg, col_reg}<20'b10011011000100011111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10011011000100011111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10011011000100100000) && ({row_reg, col_reg}<20'b10011011000101001011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10011011000101001011) && ({row_reg, col_reg}<20'b10011011000101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10011011000101001110) && ({row_reg, col_reg}<20'b10011011001101101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10011011001101101000) && ({row_reg, col_reg}<20'b10011011001101101011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10011011001101101011) && ({row_reg, col_reg}<20'b10011011001101110000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10011011001101110000) && ({row_reg, col_reg}<20'b10011011001101110011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10011011001101110011)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==20'b10011011001101110100)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10011011001101110101)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=20'b10011011001101110110) && ({row_reg, col_reg}<20'b10011011001101111111)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10011011001101111111)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10011011001110000000) && ({row_reg, col_reg}<20'b10011011010000001001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=20'b10011011010000001001) && ({row_reg, col_reg}<20'b10011011010000001011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=20'b10011011010000001011) && ({row_reg, col_reg}<20'b10011011010000001101)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10011011010000001101)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10011011010000001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10011011010000001111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=20'b10011011010000010000) && ({row_reg, col_reg}<20'b10011011010000010011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10011011010000010011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10011011010000010100) && ({row_reg, col_reg}<20'b10011011010000010111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10011011010000010111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10011011010000011000) && ({row_reg, col_reg}<20'b10011011010100011000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10011011010100011000) && ({row_reg, col_reg}<20'b10011011010100011110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10011011010100011110) && ({row_reg, col_reg}<20'b10011011010100100000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10011011010100100000) && ({row_reg, col_reg}<20'b10011011010101001010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10011011010101001010) && ({row_reg, col_reg}<20'b10011011010101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10011011010101001100) && ({row_reg, col_reg}<20'b10011011010101010000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10011011010101010000) && ({row_reg, col_reg}<20'b10011011011000110000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10011011011000110000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10011011011000110001) && ({row_reg, col_reg}<20'b10011011011000110011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10011011011000110011) && ({row_reg, col_reg}<20'b10011011011000110110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10011011011000110110) && ({row_reg, col_reg}<20'b10011011011000111000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10011011011000111000) && ({row_reg, col_reg}<20'b10011011011001101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10011011011001101000) && ({row_reg, col_reg}<20'b10011011011001101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10011011011001101100) && ({row_reg, col_reg}<20'b10011011011001101110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10011011011001101110) && ({row_reg, col_reg}<20'b10011011011101101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10011011011101101000) && ({row_reg, col_reg}<20'b10011011011101101010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10011011011101101010) && ({row_reg, col_reg}<20'b10011011011101101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10011011011101101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10011011011101101101) && ({row_reg, col_reg}<20'b10011011011101110001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10011011011101110001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==20'b10011011011101110010)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10011011011101110011)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=20'b10011011011101110100) && ({row_reg, col_reg}<20'b10011011011101111010)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=20'b10011011011101111010) && ({row_reg, col_reg}<20'b10011011011101111100)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10011011011101111100) && ({row_reg, col_reg}<20'b10011011100000001100)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=20'b10011011100000001100) && ({row_reg, col_reg}<20'b10011011100000001110)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==20'b10011011100000001110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10011011100000001111)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=20'b10011011100000010000) && ({row_reg, col_reg}<20'b10011011100000010010)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10011011100000010010) && ({row_reg, col_reg}<20'b10011011100000010100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10011011100000010100) && ({row_reg, col_reg}<20'b10011011100000010110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=20'b10011011100000010110) && ({row_reg, col_reg}<20'b10011011100000011001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10011011100000011001) && ({row_reg, col_reg}<20'b10011011100100011001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10011011100100011001) && ({row_reg, col_reg}<20'b10011011100100011111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10011011100100011111) && ({row_reg, col_reg}<20'b10011011100101001110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10011011100101001110) && ({row_reg, col_reg}<20'b10011011100101010000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10011011100101010000) && ({row_reg, col_reg}<20'b10011011101000110000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10011011101000110000) && ({row_reg, col_reg}<20'b10011011101000110011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10011011101000110011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10011011101000110100) && ({row_reg, col_reg}<20'b10011011101000110110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10011011101000110110) && ({row_reg, col_reg}<20'b10011011101001101010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10011011101001101010) && ({row_reg, col_reg}<20'b10011011101001101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10011011101001101100) && ({row_reg, col_reg}<20'b10011011101101101001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10011011101101101001) && ({row_reg, col_reg}<20'b10011011101101101011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10011011101101101011) && ({row_reg, col_reg}<20'b10011011101101101101)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=20'b10011011101101101101) && ({row_reg, col_reg}<20'b10011011101101101111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10011011101101101111) && ({row_reg, col_reg}<20'b10011011101101110001)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10011011101101110001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==20'b10011011101101110010)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=20'b10011011101101110011) && ({row_reg, col_reg}<20'b10011011101101111101)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10011011101101111101)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10011011101101111110) && ({row_reg, col_reg}<20'b10011011110000000100)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10011011110000000100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=20'b10011011110000000101) && ({row_reg, col_reg}<20'b10011011110000000111)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10011011110000000111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=20'b10011011110000001000) && ({row_reg, col_reg}<20'b10011011110000010010)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10011011110000010010)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=20'b10011011110000010011) && ({row_reg, col_reg}<20'b10011011110000010101)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==20'b10011011110000010101)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10011011110000010110) && ({row_reg, col_reg}<20'b10011011110000011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10011011110000011000) && ({row_reg, col_reg}<20'b10011011110100011110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=20'b10011011110100011110) && ({row_reg, col_reg}<20'b10011011110100100000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10011011110100100000) && ({row_reg, col_reg}<20'b10011011110101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10011011110101001101) && ({row_reg, col_reg}<20'b10011011110101010000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10011011110101010000) && ({row_reg, col_reg}<20'b10011011111000110111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==20'b10011011111000110111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10011011111000111000) && ({row_reg, col_reg}<20'b10011011111001101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10011011111001101000) && ({row_reg, col_reg}<20'b10011011111101101001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=20'b10011011111101101001) && ({row_reg, col_reg}<20'b10011011111101101011)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==20'b10011011111101101011)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10011011111101101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==20'b10011011111101101101)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=20'b10011011111101101110) && ({row_reg, col_reg}<20'b10011011111101110000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10011011111101110000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=20'b10011011111101110001) && ({row_reg, col_reg}<20'b10011011111101111111)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10011011111101111111)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10011011111110000000) && ({row_reg, col_reg}<20'b10011100000000011000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=20'b10011100000000011000) && ({row_reg, col_reg}<20'b10011100000100011110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10011100000100011110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10011100000100011111) && ({row_reg, col_reg}<20'b10011100000101001010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10011100000101001010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10011100000101001011) && ({row_reg, col_reg}<20'b10011100000101001110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10011100000101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10011100000101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10011100000101010000) && ({row_reg, col_reg}<20'b10011100001000110111)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10011100001000110111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=20'b10011100001000111000) && ({row_reg, col_reg}<20'b10011100001000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10011100001000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10011100001000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10011100001000111100) && ({row_reg, col_reg}<20'b10011100001000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10011100001000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10011100001000111111) && ({row_reg, col_reg}<20'b10011100001001100100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10011100001001100100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10011100001001100101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10011100001001100110) && ({row_reg, col_reg}<20'b10011100001001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10011100001001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10011100001001101001) && ({row_reg, col_reg}<20'b10011100001101101010)) color_data = 12'b110111011101;

		if(({row_reg, col_reg}>=20'b10011100001101101010) && ({row_reg, col_reg}<20'b10011100010100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10011100010100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10011100010100011111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10011100010100100000) && ({row_reg, col_reg}<20'b10011100010101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10011100010101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10011100010101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10011100010101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10011100010101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10011100010101010000) && ({row_reg, col_reg}<20'b10011100011000110111)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10011100011000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10011100011000111000) && ({row_reg, col_reg}<20'b10011100011000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10011100011000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10011100011000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10011100011000111100) && ({row_reg, col_reg}<20'b10011100011000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10011100011000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10011100011000111111) && ({row_reg, col_reg}<20'b10011100011001100100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10011100011001100100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10011100011001100101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10011100011001100110) && ({row_reg, col_reg}<20'b10011100011001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10011100011001101000)) color_data = 12'b101110111011;

		if(({row_reg, col_reg}>=20'b10011100011001101001) && ({row_reg, col_reg}<20'b10011100100100011001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10011100100100011001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=20'b10011100100100011010) && ({row_reg, col_reg}<20'b10011100100100011100)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10011100100100011100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==20'b10011100100100011101)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10011100100100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10011100100100011111) && ({row_reg, col_reg}<20'b10011100100101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10011100100101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10011100100101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10011100100101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10011100100101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==20'b10011100100101010000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=20'b10011100100101010001) && ({row_reg, col_reg}<20'b10011100100101010011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==20'b10011100100101010011)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10011100100101010100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=20'b10011100100101010101) && ({row_reg, col_reg}<20'b10011100100101010111)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10011100100101010111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=20'b10011100100101011000) && ({row_reg, col_reg}<20'b10011100101000110100)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10011100101000110100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=20'b10011100101000110101) && ({row_reg, col_reg}<20'b10011100101000110111)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10011100101000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10011100101000111000) && ({row_reg, col_reg}<20'b10011100101000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10011100101000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10011100101000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10011100101000111100) && ({row_reg, col_reg}<20'b10011100101000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10011100101000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10011100101000111111) && ({row_reg, col_reg}<20'b10011100101001100100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10011100101001100100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10011100101001100101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10011100101001100110) && ({row_reg, col_reg}<20'b10011100101001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10011100101001101000)) color_data = 12'b101110111011;

		if(({row_reg, col_reg}>=20'b10011100101001101001) && ({row_reg, col_reg}<20'b10011100110100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10011100110100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10011100110100011111) && ({row_reg, col_reg}<20'b10011100110101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10011100110101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10011100110101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10011100110101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10011100110101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10011100110101010000) && ({row_reg, col_reg}<20'b10011100111000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10011100111000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10011100111000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10011100111000111000) && ({row_reg, col_reg}<20'b10011100111000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10011100111000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10011100111000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10011100111000111100) && ({row_reg, col_reg}<20'b10011100111000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10011100111000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10011100111000111111) && ({row_reg, col_reg}<20'b10011100111001100100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10011100111001100100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10011100111001100101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10011100111001100110) && ({row_reg, col_reg}<20'b10011100111001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10011100111001101000)) color_data = 12'b101110111011;

		if(({row_reg, col_reg}>=20'b10011100111001101001) && ({row_reg, col_reg}<20'b10011101000100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10011101000100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10011101000100011111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10011101000100100000) && ({row_reg, col_reg}<20'b10011101000101001000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10011101000101001000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10011101000101001001) && ({row_reg, col_reg}<20'b10011101000101001110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10011101000101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10011101000101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10011101000101010000) && ({row_reg, col_reg}<20'b10011101000101010100)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10011101000101010100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=20'b10011101000101010101) && ({row_reg, col_reg}<20'b10011101001000110111)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10011101001000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10011101001000111000) && ({row_reg, col_reg}<20'b10011101001000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10011101001000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10011101001000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10011101001000111100) && ({row_reg, col_reg}<20'b10011101001000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10011101001000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10011101001000111111) && ({row_reg, col_reg}<20'b10011101001001100100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10011101001001100100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10011101001001100101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10011101001001100110) && ({row_reg, col_reg}<20'b10011101001001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10011101001001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10011101001001101001) && ({row_reg, col_reg}<20'b10011101001101101000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10011101001101101000)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10011101001101101001) && ({row_reg, col_reg}<20'b10011101010100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10011101010100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10011101010100011111) && ({row_reg, col_reg}<20'b10011101010101001000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10011101010101001000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10011101010101001001) && ({row_reg, col_reg}<20'b10011101010101001110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10011101010101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10011101010101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10011101010101010000) && ({row_reg, col_reg}<20'b10011101011000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10011101011000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10011101011000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10011101011000111000) && ({row_reg, col_reg}<20'b10011101011000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10011101011000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10011101011000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10011101011000111100) && ({row_reg, col_reg}<20'b10011101011000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10011101011000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10011101011000111111) && ({row_reg, col_reg}<20'b10011101011001100100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10011101011001100100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10011101011001100101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10011101011001100110) && ({row_reg, col_reg}<20'b10011101011001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10011101011001101000)) color_data = 12'b101110111011;

		if(({row_reg, col_reg}>=20'b10011101011001101001) && ({row_reg, col_reg}<20'b10011101100100011100)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10011101100100011100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==20'b10011101100100011101)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10011101100100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10011101100100011111) && ({row_reg, col_reg}<20'b10011101100101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10011101100101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10011101100101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10011101100101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10011101100101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10011101100101010000) && ({row_reg, col_reg}<20'b10011101100101010100)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10011101100101010100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=20'b10011101100101010101) && ({row_reg, col_reg}<20'b10011101101000110111)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10011101101000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10011101101000111000) && ({row_reg, col_reg}<20'b10011101101000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10011101101000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10011101101000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10011101101000111100) && ({row_reg, col_reg}<20'b10011101101000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10011101101000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10011101101000111111) && ({row_reg, col_reg}<20'b10011101101001100100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10011101101001100100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10011101101001100101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10011101101001100110) && ({row_reg, col_reg}<20'b10011101101001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10011101101001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10011101101001101001) && ({row_reg, col_reg}<20'b10011101101101101111)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10011101101101101111)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10011101101101110000) && ({row_reg, col_reg}<20'b10011101110100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10011101110100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10011101110100011111) && ({row_reg, col_reg}<20'b10011101110101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10011101110101001100) && ({row_reg, col_reg}<20'b10011101110101001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10011101110101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10011101110101010000) && ({row_reg, col_reg}<20'b10011101111000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10011101111000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10011101111000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10011101111000111000) && ({row_reg, col_reg}<20'b10011101111000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10011101111000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10011101111000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10011101111000111100) && ({row_reg, col_reg}<20'b10011101111000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10011101111000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10011101111000111111) && ({row_reg, col_reg}<20'b10011101111001100100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10011101111001100100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10011101111001100101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10011101111001100110) && ({row_reg, col_reg}<20'b10011101111001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10011101111001101000)) color_data = 12'b101110111011;

		if(({row_reg, col_reg}>=20'b10011101111001101001) && ({row_reg, col_reg}<20'b10011110000100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10011110000100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10011110000100011111) && ({row_reg, col_reg}<20'b10011110000101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10011110000101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10011110000101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10011110000101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10011110000101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10011110000101010000) && ({row_reg, col_reg}<20'b10011110001000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10011110001000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10011110001000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10011110001000111000) && ({row_reg, col_reg}<20'b10011110001000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10011110001000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10011110001000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10011110001000111100) && ({row_reg, col_reg}<20'b10011110001000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10011110001000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10011110001000111111) && ({row_reg, col_reg}<20'b10011110001001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10011110001001100110) && ({row_reg, col_reg}<20'b10011110001001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10011110001001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10011110001001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10011110001001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10011110001001101011) && ({row_reg, col_reg}<20'b10011110010100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10011110010100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10011110010100011111) && ({row_reg, col_reg}<20'b10011110010101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10011110010101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10011110010101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10011110010101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10011110010101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10011110010101010000) && ({row_reg, col_reg}<20'b10011110011000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10011110011000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10011110011000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10011110011000111000) && ({row_reg, col_reg}<20'b10011110011000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10011110011000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10011110011000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10011110011000111100) && ({row_reg, col_reg}<20'b10011110011000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10011110011000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10011110011000111111) && ({row_reg, col_reg}<20'b10011110011001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10011110011001100110) && ({row_reg, col_reg}<20'b10011110011001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10011110011001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10011110011001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10011110011001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10011110011001101011) && ({row_reg, col_reg}<20'b10011110100100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10011110100100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10011110100100011111) && ({row_reg, col_reg}<20'b10011110100101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10011110100101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10011110100101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10011110100101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10011110100101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10011110100101010000) && ({row_reg, col_reg}<20'b10011110101000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10011110101000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10011110101000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10011110101000111000) && ({row_reg, col_reg}<20'b10011110101000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10011110101000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10011110101000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10011110101000111100) && ({row_reg, col_reg}<20'b10011110101000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10011110101000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10011110101000111111) && ({row_reg, col_reg}<20'b10011110101001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10011110101001100110) && ({row_reg, col_reg}<20'b10011110101001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10011110101001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10011110101001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10011110101001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10011110101001101011) && ({row_reg, col_reg}<20'b10011110110100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10011110110100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10011110110100011111) && ({row_reg, col_reg}<20'b10011110110101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10011110110101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10011110110101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10011110110101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10011110110101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10011110110101010000) && ({row_reg, col_reg}<20'b10011110111000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10011110111000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10011110111000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10011110111000111000) && ({row_reg, col_reg}<20'b10011110111000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10011110111000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10011110111000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10011110111000111100) && ({row_reg, col_reg}<20'b10011110111000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10011110111000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10011110111000111111) && ({row_reg, col_reg}<20'b10011110111001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10011110111001100110) && ({row_reg, col_reg}<20'b10011110111001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10011110111001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10011110111001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10011110111001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10011110111001101011) && ({row_reg, col_reg}<20'b10011111000100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10011111000100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10011111000100011111) && ({row_reg, col_reg}<20'b10011111000101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10011111000101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10011111000101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10011111000101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10011111000101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10011111000101010000) && ({row_reg, col_reg}<20'b10011111001000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10011111001000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10011111001000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10011111001000111000) && ({row_reg, col_reg}<20'b10011111001000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10011111001000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10011111001000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10011111001000111100) && ({row_reg, col_reg}<20'b10011111001000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10011111001000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10011111001000111111) && ({row_reg, col_reg}<20'b10011111001001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10011111001001100110) && ({row_reg, col_reg}<20'b10011111001001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10011111001001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10011111001001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10011111001001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10011111001001101011) && ({row_reg, col_reg}<20'b10011111010100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10011111010100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10011111010100011111) && ({row_reg, col_reg}<20'b10011111010101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10011111010101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10011111010101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10011111010101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10011111010101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10011111010101010000) && ({row_reg, col_reg}<20'b10011111011000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10011111011000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10011111011000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10011111011000111000) && ({row_reg, col_reg}<20'b10011111011000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10011111011000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10011111011000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10011111011000111100) && ({row_reg, col_reg}<20'b10011111011000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10011111011000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10011111011000111111) && ({row_reg, col_reg}<20'b10011111011001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10011111011001100110) && ({row_reg, col_reg}<20'b10011111011001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10011111011001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10011111011001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10011111011001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10011111011001101011) && ({row_reg, col_reg}<20'b10011111100100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10011111100100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10011111100100011111) && ({row_reg, col_reg}<20'b10011111100101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10011111100101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10011111100101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10011111100101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10011111100101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10011111100101010000) && ({row_reg, col_reg}<20'b10011111101000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10011111101000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10011111101000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10011111101000111000) && ({row_reg, col_reg}<20'b10011111101000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10011111101000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10011111101000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10011111101000111100) && ({row_reg, col_reg}<20'b10011111101000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10011111101000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10011111101000111111) && ({row_reg, col_reg}<20'b10011111101001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10011111101001100110) && ({row_reg, col_reg}<20'b10011111101001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10011111101001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10011111101001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10011111101001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10011111101001101011) && ({row_reg, col_reg}<20'b10011111110100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10011111110100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10011111110100011111) && ({row_reg, col_reg}<20'b10011111110101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10011111110101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10011111110101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10011111110101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10011111110101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10011111110101010000) && ({row_reg, col_reg}<20'b10011111111000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10011111111000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10011111111000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10011111111000111000) && ({row_reg, col_reg}<20'b10011111111000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10011111111000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10011111111000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10011111111000111100) && ({row_reg, col_reg}<20'b10011111111000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10011111111000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10011111111000111111) && ({row_reg, col_reg}<20'b10011111111001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10011111111001100110) && ({row_reg, col_reg}<20'b10011111111001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10011111111001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10011111111001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10011111111001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10011111111001101011) && ({row_reg, col_reg}<20'b10100000000100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10100000000100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10100000000100011111) && ({row_reg, col_reg}<20'b10100000000101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10100000000101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10100000000101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10100000000101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10100000000101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10100000000101010000) && ({row_reg, col_reg}<20'b10100000001000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10100000001000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10100000001000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10100000001000111000) && ({row_reg, col_reg}<20'b10100000001000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10100000001000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10100000001000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10100000001000111100) && ({row_reg, col_reg}<20'b10100000001000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10100000001000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10100000001000111111) && ({row_reg, col_reg}<20'b10100000001001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10100000001001100110) && ({row_reg, col_reg}<20'b10100000001001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10100000001001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10100000001001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10100000001001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10100000001001101011) && ({row_reg, col_reg}<20'b10100000010100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10100000010100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10100000010100011111) && ({row_reg, col_reg}<20'b10100000010101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10100000010101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10100000010101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10100000010101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10100000010101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10100000010101010000) && ({row_reg, col_reg}<20'b10100000011000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10100000011000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10100000011000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10100000011000111000) && ({row_reg, col_reg}<20'b10100000011000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10100000011000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10100000011000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10100000011000111100) && ({row_reg, col_reg}<20'b10100000011000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10100000011000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10100000011000111111) && ({row_reg, col_reg}<20'b10100000011001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10100000011001100110) && ({row_reg, col_reg}<20'b10100000011001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10100000011001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10100000011001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10100000011001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10100000011001101011) && ({row_reg, col_reg}<20'b10100000100100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10100000100100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10100000100100011111) && ({row_reg, col_reg}<20'b10100000100101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10100000100101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10100000100101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10100000100101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10100000100101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10100000100101010000) && ({row_reg, col_reg}<20'b10100000101000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10100000101000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10100000101000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10100000101000111000) && ({row_reg, col_reg}<20'b10100000101000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10100000101000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10100000101000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10100000101000111100) && ({row_reg, col_reg}<20'b10100000101000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10100000101000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10100000101000111111) && ({row_reg, col_reg}<20'b10100000101001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10100000101001100110) && ({row_reg, col_reg}<20'b10100000101001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10100000101001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10100000101001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10100000101001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10100000101001101011) && ({row_reg, col_reg}<20'b10100000110100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10100000110100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10100000110100011111) && ({row_reg, col_reg}<20'b10100000110101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10100000110101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10100000110101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10100000110101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10100000110101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10100000110101010000) && ({row_reg, col_reg}<20'b10100000111000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10100000111000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10100000111000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10100000111000111000) && ({row_reg, col_reg}<20'b10100000111000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10100000111000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10100000111000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10100000111000111100) && ({row_reg, col_reg}<20'b10100000111000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10100000111000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10100000111000111111) && ({row_reg, col_reg}<20'b10100000111001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10100000111001100110) && ({row_reg, col_reg}<20'b10100000111001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10100000111001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10100000111001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10100000111001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10100000111001101011) && ({row_reg, col_reg}<20'b10100001000100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10100001000100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10100001000100011111) && ({row_reg, col_reg}<20'b10100001000101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10100001000101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10100001000101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10100001000101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10100001000101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10100001000101010000) && ({row_reg, col_reg}<20'b10100001001000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10100001001000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10100001001000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10100001001000111000) && ({row_reg, col_reg}<20'b10100001001000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10100001001000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10100001001000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10100001001000111100) && ({row_reg, col_reg}<20'b10100001001000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10100001001000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10100001001000111111) && ({row_reg, col_reg}<20'b10100001001001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10100001001001100110) && ({row_reg, col_reg}<20'b10100001001001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10100001001001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10100001001001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10100001001001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10100001001001101011) && ({row_reg, col_reg}<20'b10100001010100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10100001010100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10100001010100011111) && ({row_reg, col_reg}<20'b10100001010101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10100001010101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10100001010101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10100001010101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10100001010101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10100001010101010000) && ({row_reg, col_reg}<20'b10100001011000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10100001011000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10100001011000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10100001011000111000) && ({row_reg, col_reg}<20'b10100001011000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10100001011000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10100001011000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10100001011000111100) && ({row_reg, col_reg}<20'b10100001011000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10100001011000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10100001011000111111) && ({row_reg, col_reg}<20'b10100001011001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10100001011001100110) && ({row_reg, col_reg}<20'b10100001011001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10100001011001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10100001011001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10100001011001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10100001011001101011) && ({row_reg, col_reg}<20'b10100001100100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10100001100100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10100001100100011111) && ({row_reg, col_reg}<20'b10100001100101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10100001100101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10100001100101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10100001100101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10100001100101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10100001100101010000) && ({row_reg, col_reg}<20'b10100001101000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10100001101000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10100001101000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10100001101000111000) && ({row_reg, col_reg}<20'b10100001101000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10100001101000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10100001101000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10100001101000111100) && ({row_reg, col_reg}<20'b10100001101000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10100001101000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10100001101000111111) && ({row_reg, col_reg}<20'b10100001101001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10100001101001100110) && ({row_reg, col_reg}<20'b10100001101001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10100001101001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10100001101001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10100001101001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10100001101001101011) && ({row_reg, col_reg}<20'b10100001110100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10100001110100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10100001110100011111) && ({row_reg, col_reg}<20'b10100001110101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10100001110101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10100001110101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10100001110101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10100001110101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10100001110101010000) && ({row_reg, col_reg}<20'b10100001111000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10100001111000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10100001111000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10100001111000111000) && ({row_reg, col_reg}<20'b10100001111000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10100001111000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10100001111000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10100001111000111100) && ({row_reg, col_reg}<20'b10100001111000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10100001111000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10100001111000111111) && ({row_reg, col_reg}<20'b10100001111001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10100001111001100110) && ({row_reg, col_reg}<20'b10100001111001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10100001111001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10100001111001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10100001111001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10100001111001101011) && ({row_reg, col_reg}<20'b10100010000100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10100010000100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10100010000100011111) && ({row_reg, col_reg}<20'b10100010000101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10100010000101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10100010000101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10100010000101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10100010000101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10100010000101010000) && ({row_reg, col_reg}<20'b10100010001000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10100010001000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10100010001000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10100010001000111000) && ({row_reg, col_reg}<20'b10100010001000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10100010001000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10100010001000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10100010001000111100) && ({row_reg, col_reg}<20'b10100010001000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10100010001000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10100010001000111111) && ({row_reg, col_reg}<20'b10100010001001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10100010001001100110) && ({row_reg, col_reg}<20'b10100010001001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10100010001001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10100010001001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10100010001001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10100010001001101011) && ({row_reg, col_reg}<20'b10100010010100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10100010010100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10100010010100011111) && ({row_reg, col_reg}<20'b10100010010101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10100010010101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10100010010101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10100010010101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10100010010101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10100010010101010000) && ({row_reg, col_reg}<20'b10100010011000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10100010011000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10100010011000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10100010011000111000) && ({row_reg, col_reg}<20'b10100010011000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10100010011000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10100010011000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10100010011000111100) && ({row_reg, col_reg}<20'b10100010011000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10100010011000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10100010011000111111) && ({row_reg, col_reg}<20'b10100010011001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10100010011001100110) && ({row_reg, col_reg}<20'b10100010011001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10100010011001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10100010011001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10100010011001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10100010011001101011) && ({row_reg, col_reg}<20'b10100010100100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10100010100100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10100010100100011111) && ({row_reg, col_reg}<20'b10100010100101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10100010100101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10100010100101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10100010100101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10100010100101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10100010100101010000) && ({row_reg, col_reg}<20'b10100010101000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10100010101000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10100010101000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10100010101000111000) && ({row_reg, col_reg}<20'b10100010101000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10100010101000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10100010101000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10100010101000111100) && ({row_reg, col_reg}<20'b10100010101000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10100010101000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10100010101000111111) && ({row_reg, col_reg}<20'b10100010101001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10100010101001100110) && ({row_reg, col_reg}<20'b10100010101001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10100010101001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10100010101001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10100010101001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10100010101001101011) && ({row_reg, col_reg}<20'b10100010110100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10100010110100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10100010110100011111) && ({row_reg, col_reg}<20'b10100010110101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10100010110101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10100010110101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10100010110101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10100010110101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10100010110101010000) && ({row_reg, col_reg}<20'b10100010111000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10100010111000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10100010111000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10100010111000111000) && ({row_reg, col_reg}<20'b10100010111000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10100010111000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10100010111000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10100010111000111100) && ({row_reg, col_reg}<20'b10100010111000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10100010111000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10100010111000111111) && ({row_reg, col_reg}<20'b10100010111001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10100010111001100110) && ({row_reg, col_reg}<20'b10100010111001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10100010111001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10100010111001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10100010111001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10100010111001101011) && ({row_reg, col_reg}<20'b10100011000100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10100011000100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10100011000100011111) && ({row_reg, col_reg}<20'b10100011000101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10100011000101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10100011000101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10100011000101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10100011000101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10100011000101010000) && ({row_reg, col_reg}<20'b10100011001000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10100011001000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10100011001000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10100011001000111000) && ({row_reg, col_reg}<20'b10100011001000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10100011001000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10100011001000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10100011001000111100) && ({row_reg, col_reg}<20'b10100011001000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10100011001000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10100011001000111111) && ({row_reg, col_reg}<20'b10100011001001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10100011001001100110) && ({row_reg, col_reg}<20'b10100011001001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10100011001001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10100011001001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10100011001001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10100011001001101011) && ({row_reg, col_reg}<20'b10100011010100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10100011010100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10100011010100011111) && ({row_reg, col_reg}<20'b10100011010101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10100011010101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10100011010101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10100011010101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10100011010101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10100011010101010000) && ({row_reg, col_reg}<20'b10100011011000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10100011011000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10100011011000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10100011011000111000) && ({row_reg, col_reg}<20'b10100011011000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10100011011000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10100011011000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10100011011000111100) && ({row_reg, col_reg}<20'b10100011011000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10100011011000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10100011011000111111) && ({row_reg, col_reg}<20'b10100011011001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10100011011001100110) && ({row_reg, col_reg}<20'b10100011011001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10100011011001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10100011011001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10100011011001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10100011011001101011) && ({row_reg, col_reg}<20'b10100011100100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10100011100100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10100011100100011111) && ({row_reg, col_reg}<20'b10100011100101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10100011100101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10100011100101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10100011100101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10100011100101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10100011100101010000) && ({row_reg, col_reg}<20'b10100011101000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10100011101000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10100011101000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10100011101000111000) && ({row_reg, col_reg}<20'b10100011101000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10100011101000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10100011101000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10100011101000111100) && ({row_reg, col_reg}<20'b10100011101000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10100011101000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10100011101000111111) && ({row_reg, col_reg}<20'b10100011101001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10100011101001100110) && ({row_reg, col_reg}<20'b10100011101001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10100011101001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10100011101001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10100011101001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10100011101001101011) && ({row_reg, col_reg}<20'b10100011110100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10100011110100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10100011110100011111) && ({row_reg, col_reg}<20'b10100011110101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10100011110101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10100011110101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10100011110101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10100011110101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10100011110101010000) && ({row_reg, col_reg}<20'b10100011111000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10100011111000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10100011111000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10100011111000111000) && ({row_reg, col_reg}<20'b10100011111000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10100011111000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10100011111000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10100011111000111100) && ({row_reg, col_reg}<20'b10100011111000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10100011111000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10100011111000111111) && ({row_reg, col_reg}<20'b10100011111001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10100011111001100110) && ({row_reg, col_reg}<20'b10100011111001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10100011111001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10100011111001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10100011111001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10100011111001101011) && ({row_reg, col_reg}<20'b10100100000100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10100100000100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10100100000100011111) && ({row_reg, col_reg}<20'b10100100000101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10100100000101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10100100000101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10100100000101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10100100000101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10100100000101010000) && ({row_reg, col_reg}<20'b10100100001000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10100100001000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10100100001000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10100100001000111000) && ({row_reg, col_reg}<20'b10100100001000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10100100001000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10100100001000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10100100001000111100) && ({row_reg, col_reg}<20'b10100100001000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10100100001000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10100100001000111111) && ({row_reg, col_reg}<20'b10100100001001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10100100001001100110) && ({row_reg, col_reg}<20'b10100100001001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10100100001001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10100100001001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10100100001001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10100100001001101011) && ({row_reg, col_reg}<20'b10100100010100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10100100010100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10100100010100011111) && ({row_reg, col_reg}<20'b10100100010101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10100100010101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10100100010101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10100100010101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10100100010101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10100100010101010000) && ({row_reg, col_reg}<20'b10100100011000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10100100011000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10100100011000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10100100011000111000) && ({row_reg, col_reg}<20'b10100100011000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10100100011000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10100100011000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10100100011000111100) && ({row_reg, col_reg}<20'b10100100011000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10100100011000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10100100011000111111) && ({row_reg, col_reg}<20'b10100100011001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10100100011001100110) && ({row_reg, col_reg}<20'b10100100011001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10100100011001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10100100011001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10100100011001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10100100011001101011) && ({row_reg, col_reg}<20'b10100100100100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10100100100100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10100100100100011111) && ({row_reg, col_reg}<20'b10100100100101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10100100100101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10100100100101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10100100100101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10100100100101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10100100100101010000) && ({row_reg, col_reg}<20'b10100100101000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10100100101000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10100100101000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10100100101000111000) && ({row_reg, col_reg}<20'b10100100101000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10100100101000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10100100101000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10100100101000111100) && ({row_reg, col_reg}<20'b10100100101000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10100100101000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10100100101000111111) && ({row_reg, col_reg}<20'b10100100101001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10100100101001100110) && ({row_reg, col_reg}<20'b10100100101001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10100100101001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10100100101001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10100100101001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10100100101001101011) && ({row_reg, col_reg}<20'b10100100110100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10100100110100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10100100110100011111) && ({row_reg, col_reg}<20'b10100100110101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10100100110101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10100100110101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10100100110101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10100100110101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10100100110101010000) && ({row_reg, col_reg}<20'b10100100111000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10100100111000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10100100111000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10100100111000111000) && ({row_reg, col_reg}<20'b10100100111000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10100100111000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10100100111000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10100100111000111100) && ({row_reg, col_reg}<20'b10100100111000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10100100111000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10100100111000111111) && ({row_reg, col_reg}<20'b10100100111001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10100100111001100110) && ({row_reg, col_reg}<20'b10100100111001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10100100111001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10100100111001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10100100111001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10100100111001101011) && ({row_reg, col_reg}<20'b10100101000100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10100101000100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10100101000100011111) && ({row_reg, col_reg}<20'b10100101000101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10100101000101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10100101000101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10100101000101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10100101000101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10100101000101010000) && ({row_reg, col_reg}<20'b10100101001000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10100101001000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10100101001000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10100101001000111000) && ({row_reg, col_reg}<20'b10100101001000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10100101001000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10100101001000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10100101001000111100) && ({row_reg, col_reg}<20'b10100101001000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10100101001000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10100101001000111111) && ({row_reg, col_reg}<20'b10100101001001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10100101001001100110) && ({row_reg, col_reg}<20'b10100101001001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10100101001001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10100101001001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10100101001001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10100101001001101011) && ({row_reg, col_reg}<20'b10100101010100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10100101010100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10100101010100011111) && ({row_reg, col_reg}<20'b10100101010101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10100101010101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10100101010101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10100101010101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10100101010101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10100101010101010000) && ({row_reg, col_reg}<20'b10100101011000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10100101011000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10100101011000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10100101011000111000) && ({row_reg, col_reg}<20'b10100101011000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10100101011000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10100101011000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10100101011000111100) && ({row_reg, col_reg}<20'b10100101011000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10100101011000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10100101011000111111) && ({row_reg, col_reg}<20'b10100101011001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10100101011001100110) && ({row_reg, col_reg}<20'b10100101011001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10100101011001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10100101011001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10100101011001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10100101011001101011) && ({row_reg, col_reg}<20'b10100101100100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10100101100100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10100101100100011111) && ({row_reg, col_reg}<20'b10100101100101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10100101100101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10100101100101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10100101100101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10100101100101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10100101100101010000) && ({row_reg, col_reg}<20'b10100101101000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10100101101000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10100101101000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10100101101000111000) && ({row_reg, col_reg}<20'b10100101101000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10100101101000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10100101101000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10100101101000111100) && ({row_reg, col_reg}<20'b10100101101000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10100101101000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10100101101000111111) && ({row_reg, col_reg}<20'b10100101101001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10100101101001100110) && ({row_reg, col_reg}<20'b10100101101001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10100101101001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10100101101001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10100101101001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10100101101001101011) && ({row_reg, col_reg}<20'b10100101110100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10100101110100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10100101110100011111) && ({row_reg, col_reg}<20'b10100101110101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10100101110101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10100101110101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10100101110101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10100101110101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10100101110101010000) && ({row_reg, col_reg}<20'b10100101111000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10100101111000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10100101111000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10100101111000111000) && ({row_reg, col_reg}<20'b10100101111000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10100101111000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10100101111000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10100101111000111100) && ({row_reg, col_reg}<20'b10100101111000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10100101111000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10100101111000111111) && ({row_reg, col_reg}<20'b10100101111001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10100101111001100110) && ({row_reg, col_reg}<20'b10100101111001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10100101111001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10100101111001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10100101111001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10100101111001101011) && ({row_reg, col_reg}<20'b10100110000100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10100110000100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10100110000100011111) && ({row_reg, col_reg}<20'b10100110000101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10100110000101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10100110000101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10100110000101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10100110000101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10100110000101010000) && ({row_reg, col_reg}<20'b10100110001000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10100110001000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10100110001000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10100110001000111000) && ({row_reg, col_reg}<20'b10100110001000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10100110001000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10100110001000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10100110001000111100) && ({row_reg, col_reg}<20'b10100110001000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10100110001000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10100110001000111111) && ({row_reg, col_reg}<20'b10100110001001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10100110001001100110) && ({row_reg, col_reg}<20'b10100110001001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10100110001001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10100110001001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10100110001001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10100110001001101011) && ({row_reg, col_reg}<20'b10100110010100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10100110010100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10100110010100011111) && ({row_reg, col_reg}<20'b10100110010101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10100110010101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10100110010101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10100110010101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10100110010101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10100110010101010000) && ({row_reg, col_reg}<20'b10100110011000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10100110011000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10100110011000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10100110011000111000) && ({row_reg, col_reg}<20'b10100110011000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10100110011000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10100110011000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10100110011000111100) && ({row_reg, col_reg}<20'b10100110011000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10100110011000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10100110011000111111) && ({row_reg, col_reg}<20'b10100110011001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10100110011001100110) && ({row_reg, col_reg}<20'b10100110011001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10100110011001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10100110011001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10100110011001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10100110011001101011) && ({row_reg, col_reg}<20'b10100110100100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10100110100100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10100110100100011111) && ({row_reg, col_reg}<20'b10100110100101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10100110100101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10100110100101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10100110100101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10100110100101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10100110100101010000) && ({row_reg, col_reg}<20'b10100110101000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10100110101000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10100110101000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10100110101000111000) && ({row_reg, col_reg}<20'b10100110101000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10100110101000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10100110101000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10100110101000111100) && ({row_reg, col_reg}<20'b10100110101000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10100110101000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10100110101000111111) && ({row_reg, col_reg}<20'b10100110101001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10100110101001100110) && ({row_reg, col_reg}<20'b10100110101001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10100110101001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10100110101001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10100110101001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10100110101001101011) && ({row_reg, col_reg}<20'b10100110110100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10100110110100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10100110110100011111) && ({row_reg, col_reg}<20'b10100110110101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10100110110101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10100110110101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10100110110101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10100110110101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10100110110101010000) && ({row_reg, col_reg}<20'b10100110111000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10100110111000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10100110111000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10100110111000111000) && ({row_reg, col_reg}<20'b10100110111000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10100110111000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10100110111000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10100110111000111100) && ({row_reg, col_reg}<20'b10100110111000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10100110111000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10100110111000111111) && ({row_reg, col_reg}<20'b10100110111001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10100110111001100110) && ({row_reg, col_reg}<20'b10100110111001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10100110111001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10100110111001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10100110111001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10100110111001101011) && ({row_reg, col_reg}<20'b10100111000100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10100111000100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10100111000100011111) && ({row_reg, col_reg}<20'b10100111000101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10100111000101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10100111000101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10100111000101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10100111000101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10100111000101010000) && ({row_reg, col_reg}<20'b10100111001000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10100111001000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10100111001000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10100111001000111000) && ({row_reg, col_reg}<20'b10100111001000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10100111001000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10100111001000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10100111001000111100) && ({row_reg, col_reg}<20'b10100111001000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10100111001000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10100111001000111111) && ({row_reg, col_reg}<20'b10100111001001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10100111001001100110) && ({row_reg, col_reg}<20'b10100111001001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10100111001001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10100111001001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10100111001001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10100111001001101011) && ({row_reg, col_reg}<20'b10100111010100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10100111010100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10100111010100011111) && ({row_reg, col_reg}<20'b10100111010101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10100111010101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10100111010101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10100111010101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10100111010101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10100111010101010000) && ({row_reg, col_reg}<20'b10100111011000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10100111011000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10100111011000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10100111011000111000) && ({row_reg, col_reg}<20'b10100111011000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10100111011000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10100111011000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10100111011000111100) && ({row_reg, col_reg}<20'b10100111011000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10100111011000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10100111011000111111) && ({row_reg, col_reg}<20'b10100111011001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10100111011001100110) && ({row_reg, col_reg}<20'b10100111011001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10100111011001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10100111011001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10100111011001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10100111011001101011) && ({row_reg, col_reg}<20'b10100111100100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10100111100100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10100111100100011111) && ({row_reg, col_reg}<20'b10100111100101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10100111100101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10100111100101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10100111100101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10100111100101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10100111100101010000) && ({row_reg, col_reg}<20'b10100111101000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10100111101000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10100111101000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10100111101000111000) && ({row_reg, col_reg}<20'b10100111101000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10100111101000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10100111101000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10100111101000111100) && ({row_reg, col_reg}<20'b10100111101000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10100111101000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10100111101000111111) && ({row_reg, col_reg}<20'b10100111101001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10100111101001100110) && ({row_reg, col_reg}<20'b10100111101001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10100111101001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10100111101001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10100111101001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10100111101001101011) && ({row_reg, col_reg}<20'b10100111110100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10100111110100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10100111110100011111) && ({row_reg, col_reg}<20'b10100111110101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10100111110101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10100111110101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10100111110101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10100111110101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10100111110101010000) && ({row_reg, col_reg}<20'b10100111111000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10100111111000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10100111111000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10100111111000111000) && ({row_reg, col_reg}<20'b10100111111000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10100111111000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10100111111000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10100111111000111100) && ({row_reg, col_reg}<20'b10100111111000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10100111111000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10100111111000111111) && ({row_reg, col_reg}<20'b10100111111001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10100111111001100110) && ({row_reg, col_reg}<20'b10100111111001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10100111111001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10100111111001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10100111111001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10100111111001101011) && ({row_reg, col_reg}<20'b10101000000100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10101000000100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10101000000100011111) && ({row_reg, col_reg}<20'b10101000000101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10101000000101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10101000000101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10101000000101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10101000000101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10101000000101010000) && ({row_reg, col_reg}<20'b10101000001000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10101000001000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10101000001000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10101000001000111000) && ({row_reg, col_reg}<20'b10101000001000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10101000001000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10101000001000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10101000001000111100) && ({row_reg, col_reg}<20'b10101000001000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10101000001000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10101000001000111111) && ({row_reg, col_reg}<20'b10101000001001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10101000001001100110) && ({row_reg, col_reg}<20'b10101000001001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10101000001001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10101000001001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10101000001001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10101000001001101011) && ({row_reg, col_reg}<20'b10101000010100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10101000010100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10101000010100011111) && ({row_reg, col_reg}<20'b10101000010101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10101000010101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10101000010101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10101000010101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10101000010101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10101000010101010000) && ({row_reg, col_reg}<20'b10101000011000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10101000011000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10101000011000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10101000011000111000) && ({row_reg, col_reg}<20'b10101000011000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10101000011000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10101000011000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10101000011000111100) && ({row_reg, col_reg}<20'b10101000011000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10101000011000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10101000011000111111) && ({row_reg, col_reg}<20'b10101000011001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10101000011001100110) && ({row_reg, col_reg}<20'b10101000011001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10101000011001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10101000011001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10101000011001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10101000011001101011) && ({row_reg, col_reg}<20'b10101000100100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10101000100100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10101000100100011111) && ({row_reg, col_reg}<20'b10101000100101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10101000100101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10101000100101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10101000100101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10101000100101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10101000100101010000) && ({row_reg, col_reg}<20'b10101000101000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10101000101000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10101000101000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10101000101000111000) && ({row_reg, col_reg}<20'b10101000101000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10101000101000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10101000101000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10101000101000111100) && ({row_reg, col_reg}<20'b10101000101000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10101000101000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10101000101000111111) && ({row_reg, col_reg}<20'b10101000101001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10101000101001100110) && ({row_reg, col_reg}<20'b10101000101001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10101000101001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10101000101001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10101000101001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10101000101001101011) && ({row_reg, col_reg}<20'b10101000110100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10101000110100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10101000110100011111) && ({row_reg, col_reg}<20'b10101000110101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10101000110101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10101000110101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10101000110101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10101000110101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10101000110101010000) && ({row_reg, col_reg}<20'b10101000111000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10101000111000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10101000111000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10101000111000111000) && ({row_reg, col_reg}<20'b10101000111000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10101000111000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10101000111000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10101000111000111100) && ({row_reg, col_reg}<20'b10101000111000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10101000111000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10101000111000111111) && ({row_reg, col_reg}<20'b10101000111001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10101000111001100110) && ({row_reg, col_reg}<20'b10101000111001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10101000111001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10101000111001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10101000111001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10101000111001101011) && ({row_reg, col_reg}<20'b10101001000100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10101001000100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10101001000100011111) && ({row_reg, col_reg}<20'b10101001000101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10101001000101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10101001000101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10101001000101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10101001000101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10101001000101010000) && ({row_reg, col_reg}<20'b10101001001000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10101001001000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10101001001000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10101001001000111000) && ({row_reg, col_reg}<20'b10101001001000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10101001001000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10101001001000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10101001001000111100) && ({row_reg, col_reg}<20'b10101001001000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10101001001000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10101001001000111111) && ({row_reg, col_reg}<20'b10101001001001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10101001001001100110) && ({row_reg, col_reg}<20'b10101001001001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10101001001001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10101001001001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10101001001001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10101001001001101011) && ({row_reg, col_reg}<20'b10101001010100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10101001010100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10101001010100011111) && ({row_reg, col_reg}<20'b10101001010101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10101001010101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10101001010101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10101001010101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10101001010101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10101001010101010000) && ({row_reg, col_reg}<20'b10101001011000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10101001011000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10101001011000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10101001011000111000) && ({row_reg, col_reg}<20'b10101001011000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10101001011000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10101001011000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10101001011000111100) && ({row_reg, col_reg}<20'b10101001011000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10101001011000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10101001011000111111) && ({row_reg, col_reg}<20'b10101001011001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10101001011001100110) && ({row_reg, col_reg}<20'b10101001011001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10101001011001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10101001011001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10101001011001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10101001011001101011) && ({row_reg, col_reg}<20'b10101001100100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10101001100100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10101001100100011111) && ({row_reg, col_reg}<20'b10101001100101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10101001100101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10101001100101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10101001100101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10101001100101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10101001100101010000) && ({row_reg, col_reg}<20'b10101001101000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10101001101000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10101001101000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10101001101000111000) && ({row_reg, col_reg}<20'b10101001101000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10101001101000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10101001101000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10101001101000111100) && ({row_reg, col_reg}<20'b10101001101000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10101001101000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10101001101000111111) && ({row_reg, col_reg}<20'b10101001101001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10101001101001100110) && ({row_reg, col_reg}<20'b10101001101001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10101001101001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10101001101001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10101001101001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10101001101001101011) && ({row_reg, col_reg}<20'b10101001110100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10101001110100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10101001110100011111) && ({row_reg, col_reg}<20'b10101001110101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10101001110101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10101001110101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10101001110101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10101001110101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10101001110101010000) && ({row_reg, col_reg}<20'b10101001111000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10101001111000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10101001111000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10101001111000111000) && ({row_reg, col_reg}<20'b10101001111000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10101001111000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10101001111000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10101001111000111100) && ({row_reg, col_reg}<20'b10101001111000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10101001111000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10101001111000111111) && ({row_reg, col_reg}<20'b10101001111001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10101001111001100110) && ({row_reg, col_reg}<20'b10101001111001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10101001111001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10101001111001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10101001111001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10101001111001101011) && ({row_reg, col_reg}<20'b10101010000100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10101010000100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10101010000100011111) && ({row_reg, col_reg}<20'b10101010000101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10101010000101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10101010000101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10101010000101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10101010000101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10101010000101010000) && ({row_reg, col_reg}<20'b10101010001000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10101010001000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10101010001000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10101010001000111000) && ({row_reg, col_reg}<20'b10101010001000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10101010001000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10101010001000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10101010001000111100) && ({row_reg, col_reg}<20'b10101010001000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10101010001000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10101010001000111111) && ({row_reg, col_reg}<20'b10101010001001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10101010001001100110) && ({row_reg, col_reg}<20'b10101010001001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10101010001001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10101010001001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10101010001001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10101010001001101011) && ({row_reg, col_reg}<20'b10101010010100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10101010010100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10101010010100011111) && ({row_reg, col_reg}<20'b10101010010101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10101010010101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10101010010101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10101010010101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10101010010101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10101010010101010000) && ({row_reg, col_reg}<20'b10101010011000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10101010011000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10101010011000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10101010011000111000) && ({row_reg, col_reg}<20'b10101010011000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10101010011000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10101010011000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10101010011000111100) && ({row_reg, col_reg}<20'b10101010011000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10101010011000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10101010011000111111) && ({row_reg, col_reg}<20'b10101010011001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10101010011001100110) && ({row_reg, col_reg}<20'b10101010011001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10101010011001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10101010011001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10101010011001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10101010011001101011) && ({row_reg, col_reg}<20'b10101010100100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10101010100100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10101010100100011111) && ({row_reg, col_reg}<20'b10101010100101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10101010100101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10101010100101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10101010100101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10101010100101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10101010100101010000) && ({row_reg, col_reg}<20'b10101010101000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10101010101000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10101010101000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10101010101000111000) && ({row_reg, col_reg}<20'b10101010101000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10101010101000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10101010101000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10101010101000111100) && ({row_reg, col_reg}<20'b10101010101000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10101010101000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10101010101000111111) && ({row_reg, col_reg}<20'b10101010101001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10101010101001100110) && ({row_reg, col_reg}<20'b10101010101001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10101010101001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10101010101001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10101010101001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10101010101001101011) && ({row_reg, col_reg}<20'b10101010110100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10101010110100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10101010110100011111) && ({row_reg, col_reg}<20'b10101010110101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10101010110101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10101010110101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10101010110101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10101010110101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10101010110101010000) && ({row_reg, col_reg}<20'b10101010111000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10101010111000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10101010111000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10101010111000111000) && ({row_reg, col_reg}<20'b10101010111000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10101010111000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10101010111000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10101010111000111100) && ({row_reg, col_reg}<20'b10101010111000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10101010111000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10101010111000111111) && ({row_reg, col_reg}<20'b10101010111001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10101010111001100110) && ({row_reg, col_reg}<20'b10101010111001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10101010111001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10101010111001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10101010111001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10101010111001101011) && ({row_reg, col_reg}<20'b10101011000100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10101011000100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10101011000100011111) && ({row_reg, col_reg}<20'b10101011000101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10101011000101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10101011000101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10101011000101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10101011000101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10101011000101010000) && ({row_reg, col_reg}<20'b10101011001000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10101011001000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10101011001000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10101011001000111000) && ({row_reg, col_reg}<20'b10101011001000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10101011001000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10101011001000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10101011001000111100) && ({row_reg, col_reg}<20'b10101011001000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10101011001000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10101011001000111111) && ({row_reg, col_reg}<20'b10101011001001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10101011001001100110) && ({row_reg, col_reg}<20'b10101011001001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10101011001001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10101011001001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10101011001001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10101011001001101011) && ({row_reg, col_reg}<20'b10101011010100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10101011010100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10101011010100011111) && ({row_reg, col_reg}<20'b10101011010101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10101011010101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10101011010101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10101011010101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10101011010101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10101011010101010000) && ({row_reg, col_reg}<20'b10101011011000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10101011011000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10101011011000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10101011011000111000) && ({row_reg, col_reg}<20'b10101011011000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10101011011000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10101011011000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10101011011000111100) && ({row_reg, col_reg}<20'b10101011011000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10101011011000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10101011011000111111) && ({row_reg, col_reg}<20'b10101011011001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10101011011001100110) && ({row_reg, col_reg}<20'b10101011011001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10101011011001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10101011011001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10101011011001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10101011011001101011) && ({row_reg, col_reg}<20'b10101011100100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10101011100100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10101011100100011111) && ({row_reg, col_reg}<20'b10101011100101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10101011100101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10101011100101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10101011100101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10101011100101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10101011100101010000) && ({row_reg, col_reg}<20'b10101011101000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10101011101000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10101011101000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10101011101000111000) && ({row_reg, col_reg}<20'b10101011101000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10101011101000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10101011101000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10101011101000111100) && ({row_reg, col_reg}<20'b10101011101000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10101011101000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10101011101000111111) && ({row_reg, col_reg}<20'b10101011101001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10101011101001100110) && ({row_reg, col_reg}<20'b10101011101001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10101011101001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10101011101001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10101011101001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10101011101001101011) && ({row_reg, col_reg}<20'b10101011110100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10101011110100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10101011110100011111) && ({row_reg, col_reg}<20'b10101011110101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10101011110101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10101011110101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10101011110101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10101011110101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10101011110101010000) && ({row_reg, col_reg}<20'b10101011111000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10101011111000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10101011111000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10101011111000111000) && ({row_reg, col_reg}<20'b10101011111000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10101011111000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10101011111000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10101011111000111100) && ({row_reg, col_reg}<20'b10101011111000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10101011111000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10101011111000111111) && ({row_reg, col_reg}<20'b10101011111001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10101011111001100110) && ({row_reg, col_reg}<20'b10101011111001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10101011111001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10101011111001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10101011111001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10101011111001101011) && ({row_reg, col_reg}<20'b10101100000100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10101100000100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10101100000100011111) && ({row_reg, col_reg}<20'b10101100000101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10101100000101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10101100000101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10101100000101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10101100000101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10101100000101010000) && ({row_reg, col_reg}<20'b10101100001000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10101100001000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10101100001000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10101100001000111000) && ({row_reg, col_reg}<20'b10101100001000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10101100001000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10101100001000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10101100001000111100) && ({row_reg, col_reg}<20'b10101100001000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10101100001000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10101100001000111111) && ({row_reg, col_reg}<20'b10101100001001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10101100001001100110) && ({row_reg, col_reg}<20'b10101100001001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10101100001001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10101100001001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10101100001001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10101100001001101011) && ({row_reg, col_reg}<20'b10101100010100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10101100010100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10101100010100011111) && ({row_reg, col_reg}<20'b10101100010101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10101100010101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10101100010101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10101100010101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10101100010101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10101100010101010000) && ({row_reg, col_reg}<20'b10101100011000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10101100011000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10101100011000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10101100011000111000) && ({row_reg, col_reg}<20'b10101100011000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10101100011000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10101100011000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10101100011000111100) && ({row_reg, col_reg}<20'b10101100011000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10101100011000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10101100011000111111) && ({row_reg, col_reg}<20'b10101100011001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10101100011001100110) && ({row_reg, col_reg}<20'b10101100011001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10101100011001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10101100011001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10101100011001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10101100011001101011) && ({row_reg, col_reg}<20'b10101100100100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10101100100100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10101100100100011111) && ({row_reg, col_reg}<20'b10101100100101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10101100100101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10101100100101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10101100100101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10101100100101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10101100100101010000) && ({row_reg, col_reg}<20'b10101100101000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10101100101000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10101100101000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10101100101000111000) && ({row_reg, col_reg}<20'b10101100101000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10101100101000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10101100101000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10101100101000111100) && ({row_reg, col_reg}<20'b10101100101000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10101100101000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10101100101000111111) && ({row_reg, col_reg}<20'b10101100101001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10101100101001100110) && ({row_reg, col_reg}<20'b10101100101001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10101100101001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10101100101001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10101100101001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10101100101001101011) && ({row_reg, col_reg}<20'b10101100110100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10101100110100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10101100110100011111) && ({row_reg, col_reg}<20'b10101100110101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10101100110101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10101100110101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10101100110101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10101100110101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10101100110101010000) && ({row_reg, col_reg}<20'b10101100111000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10101100111000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10101100111000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10101100111000111000) && ({row_reg, col_reg}<20'b10101100111000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10101100111000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10101100111000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10101100111000111100) && ({row_reg, col_reg}<20'b10101100111000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10101100111000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10101100111000111111) && ({row_reg, col_reg}<20'b10101100111001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10101100111001100110) && ({row_reg, col_reg}<20'b10101100111001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10101100111001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10101100111001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10101100111001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10101100111001101011) && ({row_reg, col_reg}<20'b10101101000100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10101101000100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10101101000100011111) && ({row_reg, col_reg}<20'b10101101000101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10101101000101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10101101000101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10101101000101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10101101000101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10101101000101010000) && ({row_reg, col_reg}<20'b10101101001000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10101101001000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10101101001000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10101101001000111000) && ({row_reg, col_reg}<20'b10101101001000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10101101001000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10101101001000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10101101001000111100) && ({row_reg, col_reg}<20'b10101101001000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10101101001000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10101101001000111111) && ({row_reg, col_reg}<20'b10101101001001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10101101001001100110) && ({row_reg, col_reg}<20'b10101101001001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10101101001001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10101101001001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10101101001001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10101101001001101011) && ({row_reg, col_reg}<20'b10101101010100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10101101010100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10101101010100011111) && ({row_reg, col_reg}<20'b10101101010101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10101101010101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10101101010101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10101101010101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10101101010101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10101101010101010000) && ({row_reg, col_reg}<20'b10101101011000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10101101011000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10101101011000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10101101011000111000) && ({row_reg, col_reg}<20'b10101101011000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10101101011000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10101101011000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10101101011000111100) && ({row_reg, col_reg}<20'b10101101011000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10101101011000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10101101011000111111) && ({row_reg, col_reg}<20'b10101101011001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10101101011001100110) && ({row_reg, col_reg}<20'b10101101011001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10101101011001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10101101011001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10101101011001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10101101011001101011) && ({row_reg, col_reg}<20'b10101101100100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10101101100100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10101101100100011111) && ({row_reg, col_reg}<20'b10101101100101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10101101100101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10101101100101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10101101100101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10101101100101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10101101100101010000) && ({row_reg, col_reg}<20'b10101101101000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10101101101000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10101101101000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10101101101000111000) && ({row_reg, col_reg}<20'b10101101101000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10101101101000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10101101101000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10101101101000111100) && ({row_reg, col_reg}<20'b10101101101000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10101101101000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10101101101000111111) && ({row_reg, col_reg}<20'b10101101101001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10101101101001100110) && ({row_reg, col_reg}<20'b10101101101001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10101101101001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10101101101001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10101101101001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10101101101001101011) && ({row_reg, col_reg}<20'b10101101110100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10101101110100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10101101110100011111) && ({row_reg, col_reg}<20'b10101101110101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10101101110101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10101101110101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10101101110101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10101101110101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10101101110101010000) && ({row_reg, col_reg}<20'b10101101111000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10101101111000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10101101111000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10101101111000111000) && ({row_reg, col_reg}<20'b10101101111000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10101101111000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10101101111000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10101101111000111100) && ({row_reg, col_reg}<20'b10101101111000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10101101111000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10101101111000111111) && ({row_reg, col_reg}<20'b10101101111001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10101101111001100110) && ({row_reg, col_reg}<20'b10101101111001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10101101111001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10101101111001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10101101111001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10101101111001101011) && ({row_reg, col_reg}<20'b10101110000100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10101110000100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10101110000100011111) && ({row_reg, col_reg}<20'b10101110000101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10101110000101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10101110000101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10101110000101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10101110000101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10101110000101010000) && ({row_reg, col_reg}<20'b10101110001000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10101110001000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10101110001000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10101110001000111000) && ({row_reg, col_reg}<20'b10101110001000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10101110001000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10101110001000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10101110001000111100) && ({row_reg, col_reg}<20'b10101110001000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10101110001000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10101110001000111111) && ({row_reg, col_reg}<20'b10101110001001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10101110001001100110) && ({row_reg, col_reg}<20'b10101110001001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10101110001001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10101110001001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10101110001001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10101110001001101011) && ({row_reg, col_reg}<20'b10101110010100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10101110010100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10101110010100011111) && ({row_reg, col_reg}<20'b10101110010101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10101110010101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10101110010101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10101110010101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10101110010101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10101110010101010000) && ({row_reg, col_reg}<20'b10101110011000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10101110011000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10101110011000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10101110011000111000) && ({row_reg, col_reg}<20'b10101110011000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10101110011000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10101110011000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10101110011000111100) && ({row_reg, col_reg}<20'b10101110011000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10101110011000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10101110011000111111) && ({row_reg, col_reg}<20'b10101110011001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10101110011001100110) && ({row_reg, col_reg}<20'b10101110011001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10101110011001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10101110011001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10101110011001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10101110011001101011) && ({row_reg, col_reg}<20'b10101110100100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10101110100100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10101110100100011111) && ({row_reg, col_reg}<20'b10101110100101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10101110100101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10101110100101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10101110100101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10101110100101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10101110100101010000) && ({row_reg, col_reg}<20'b10101110101000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10101110101000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10101110101000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10101110101000111000) && ({row_reg, col_reg}<20'b10101110101000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10101110101000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10101110101000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10101110101000111100) && ({row_reg, col_reg}<20'b10101110101000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10101110101000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10101110101000111111) && ({row_reg, col_reg}<20'b10101110101001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10101110101001100110) && ({row_reg, col_reg}<20'b10101110101001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10101110101001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10101110101001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10101110101001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10101110101001101011) && ({row_reg, col_reg}<20'b10101110110100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10101110110100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10101110110100011111) && ({row_reg, col_reg}<20'b10101110110101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10101110110101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10101110110101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10101110110101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10101110110101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10101110110101010000) && ({row_reg, col_reg}<20'b10101110111000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10101110111000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10101110111000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10101110111000111000) && ({row_reg, col_reg}<20'b10101110111000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10101110111000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10101110111000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10101110111000111100) && ({row_reg, col_reg}<20'b10101110111000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10101110111000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10101110111000111111) && ({row_reg, col_reg}<20'b10101110111001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10101110111001100110) && ({row_reg, col_reg}<20'b10101110111001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10101110111001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10101110111001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10101110111001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10101110111001101011) && ({row_reg, col_reg}<20'b10101111000100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10101111000100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10101111000100011111) && ({row_reg, col_reg}<20'b10101111000101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10101111000101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10101111000101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10101111000101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10101111000101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10101111000101010000) && ({row_reg, col_reg}<20'b10101111001000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10101111001000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10101111001000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10101111001000111000) && ({row_reg, col_reg}<20'b10101111001000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10101111001000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10101111001000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10101111001000111100) && ({row_reg, col_reg}<20'b10101111001000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10101111001000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10101111001000111111) && ({row_reg, col_reg}<20'b10101111001001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10101111001001100110) && ({row_reg, col_reg}<20'b10101111001001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10101111001001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10101111001001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10101111001001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10101111001001101011) && ({row_reg, col_reg}<20'b10101111010100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10101111010100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10101111010100011111) && ({row_reg, col_reg}<20'b10101111010101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10101111010101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10101111010101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10101111010101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10101111010101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10101111010101010000) && ({row_reg, col_reg}<20'b10101111011000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10101111011000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10101111011000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10101111011000111000) && ({row_reg, col_reg}<20'b10101111011000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10101111011000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10101111011000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10101111011000111100) && ({row_reg, col_reg}<20'b10101111011000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10101111011000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10101111011000111111) && ({row_reg, col_reg}<20'b10101111011001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10101111011001100110) && ({row_reg, col_reg}<20'b10101111011001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10101111011001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10101111011001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10101111011001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10101111011001101011) && ({row_reg, col_reg}<20'b10101111100100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10101111100100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10101111100100011111) && ({row_reg, col_reg}<20'b10101111100101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10101111100101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10101111100101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10101111100101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10101111100101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10101111100101010000) && ({row_reg, col_reg}<20'b10101111101000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10101111101000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10101111101000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10101111101000111000) && ({row_reg, col_reg}<20'b10101111101000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10101111101000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10101111101000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10101111101000111100) && ({row_reg, col_reg}<20'b10101111101000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10101111101000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10101111101000111111) && ({row_reg, col_reg}<20'b10101111101001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10101111101001100110) && ({row_reg, col_reg}<20'b10101111101001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10101111101001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10101111101001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10101111101001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10101111101001101011) && ({row_reg, col_reg}<20'b10101111110100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10101111110100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10101111110100011111) && ({row_reg, col_reg}<20'b10101111110101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10101111110101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10101111110101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10101111110101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10101111110101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10101111110101010000) && ({row_reg, col_reg}<20'b10101111111000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10101111111000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10101111111000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10101111111000111000) && ({row_reg, col_reg}<20'b10101111111000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10101111111000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10101111111000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10101111111000111100) && ({row_reg, col_reg}<20'b10101111111000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10101111111000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10101111111000111111) && ({row_reg, col_reg}<20'b10101111111001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10101111111001100110) && ({row_reg, col_reg}<20'b10101111111001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10101111111001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10101111111001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10101111111001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10101111111001101011) && ({row_reg, col_reg}<20'b10110000000100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10110000000100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10110000000100011111) && ({row_reg, col_reg}<20'b10110000000101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10110000000101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10110000000101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10110000000101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10110000000101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10110000000101010000) && ({row_reg, col_reg}<20'b10110000001000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10110000001000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10110000001000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10110000001000111000) && ({row_reg, col_reg}<20'b10110000001000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10110000001000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10110000001000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10110000001000111100) && ({row_reg, col_reg}<20'b10110000001000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10110000001000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10110000001000111111) && ({row_reg, col_reg}<20'b10110000001001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10110000001001100110) && ({row_reg, col_reg}<20'b10110000001001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10110000001001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10110000001001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10110000001001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10110000001001101011) && ({row_reg, col_reg}<20'b10110000010100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10110000010100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10110000010100011111) && ({row_reg, col_reg}<20'b10110000010101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10110000010101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10110000010101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10110000010101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10110000010101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10110000010101010000) && ({row_reg, col_reg}<20'b10110000011000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10110000011000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10110000011000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10110000011000111000) && ({row_reg, col_reg}<20'b10110000011000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10110000011000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10110000011000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10110000011000111100) && ({row_reg, col_reg}<20'b10110000011000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10110000011000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10110000011000111111) && ({row_reg, col_reg}<20'b10110000011001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10110000011001100110) && ({row_reg, col_reg}<20'b10110000011001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10110000011001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10110000011001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10110000011001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10110000011001101011) && ({row_reg, col_reg}<20'b10110000100100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10110000100100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10110000100100011111) && ({row_reg, col_reg}<20'b10110000100101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10110000100101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10110000100101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10110000100101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10110000100101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10110000100101010000) && ({row_reg, col_reg}<20'b10110000101000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10110000101000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10110000101000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10110000101000111000) && ({row_reg, col_reg}<20'b10110000101000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10110000101000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10110000101000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10110000101000111100) && ({row_reg, col_reg}<20'b10110000101000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10110000101000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10110000101000111111) && ({row_reg, col_reg}<20'b10110000101001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10110000101001100110) && ({row_reg, col_reg}<20'b10110000101001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10110000101001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10110000101001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10110000101001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10110000101001101011) && ({row_reg, col_reg}<20'b10110000110100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10110000110100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10110000110100011111) && ({row_reg, col_reg}<20'b10110000110101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10110000110101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10110000110101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10110000110101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10110000110101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10110000110101010000) && ({row_reg, col_reg}<20'b10110000111000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10110000111000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10110000111000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10110000111000111000) && ({row_reg, col_reg}<20'b10110000111000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10110000111000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10110000111000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10110000111000111100) && ({row_reg, col_reg}<20'b10110000111000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10110000111000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10110000111000111111) && ({row_reg, col_reg}<20'b10110000111001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10110000111001100110) && ({row_reg, col_reg}<20'b10110000111001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10110000111001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10110000111001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10110000111001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10110000111001101011) && ({row_reg, col_reg}<20'b10110001000100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10110001000100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10110001000100011111) && ({row_reg, col_reg}<20'b10110001000101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10110001000101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10110001000101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10110001000101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10110001000101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10110001000101010000) && ({row_reg, col_reg}<20'b10110001001000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10110001001000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10110001001000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10110001001000111000) && ({row_reg, col_reg}<20'b10110001001000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10110001001000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10110001001000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10110001001000111100) && ({row_reg, col_reg}<20'b10110001001000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10110001001000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10110001001000111111) && ({row_reg, col_reg}<20'b10110001001001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10110001001001100110) && ({row_reg, col_reg}<20'b10110001001001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10110001001001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10110001001001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10110001001001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10110001001001101011) && ({row_reg, col_reg}<20'b10110001010100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10110001010100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10110001010100011111) && ({row_reg, col_reg}<20'b10110001010101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10110001010101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10110001010101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10110001010101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10110001010101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10110001010101010000) && ({row_reg, col_reg}<20'b10110001011000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10110001011000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10110001011000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10110001011000111000) && ({row_reg, col_reg}<20'b10110001011000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10110001011000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10110001011000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10110001011000111100) && ({row_reg, col_reg}<20'b10110001011000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10110001011000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10110001011000111111) && ({row_reg, col_reg}<20'b10110001011001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10110001011001100110) && ({row_reg, col_reg}<20'b10110001011001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10110001011001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10110001011001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10110001011001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10110001011001101011) && ({row_reg, col_reg}<20'b10110001100100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10110001100100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10110001100100011111) && ({row_reg, col_reg}<20'b10110001100101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10110001100101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10110001100101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10110001100101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10110001100101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10110001100101010000) && ({row_reg, col_reg}<20'b10110001101000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10110001101000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10110001101000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10110001101000111000) && ({row_reg, col_reg}<20'b10110001101000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10110001101000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10110001101000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10110001101000111100) && ({row_reg, col_reg}<20'b10110001101000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10110001101000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10110001101000111111) && ({row_reg, col_reg}<20'b10110001101001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10110001101001100110) && ({row_reg, col_reg}<20'b10110001101001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10110001101001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10110001101001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10110001101001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10110001101001101011) && ({row_reg, col_reg}<20'b10110001110100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10110001110100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10110001110100011111) && ({row_reg, col_reg}<20'b10110001110101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10110001110101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10110001110101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10110001110101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10110001110101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10110001110101010000) && ({row_reg, col_reg}<20'b10110001111000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10110001111000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10110001111000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10110001111000111000) && ({row_reg, col_reg}<20'b10110001111000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10110001111000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10110001111000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10110001111000111100) && ({row_reg, col_reg}<20'b10110001111000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10110001111000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10110001111000111111) && ({row_reg, col_reg}<20'b10110001111001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10110001111001100110) && ({row_reg, col_reg}<20'b10110001111001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10110001111001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10110001111001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10110001111001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10110001111001101011) && ({row_reg, col_reg}<20'b10110010000100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10110010000100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10110010000100011111) && ({row_reg, col_reg}<20'b10110010000101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10110010000101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10110010000101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10110010000101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10110010000101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10110010000101010000) && ({row_reg, col_reg}<20'b10110010001000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10110010001000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10110010001000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10110010001000111000) && ({row_reg, col_reg}<20'b10110010001000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10110010001000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10110010001000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10110010001000111100) && ({row_reg, col_reg}<20'b10110010001000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10110010001000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10110010001000111111) && ({row_reg, col_reg}<20'b10110010001001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10110010001001100110) && ({row_reg, col_reg}<20'b10110010001001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10110010001001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10110010001001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10110010001001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10110010001001101011) && ({row_reg, col_reg}<20'b10110010010100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10110010010100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10110010010100011111) && ({row_reg, col_reg}<20'b10110010010101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10110010010101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10110010010101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10110010010101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10110010010101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10110010010101010000) && ({row_reg, col_reg}<20'b10110010011000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10110010011000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10110010011000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10110010011000111000) && ({row_reg, col_reg}<20'b10110010011000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10110010011000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10110010011000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10110010011000111100) && ({row_reg, col_reg}<20'b10110010011000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10110010011000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10110010011000111111) && ({row_reg, col_reg}<20'b10110010011001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10110010011001100110) && ({row_reg, col_reg}<20'b10110010011001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10110010011001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10110010011001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10110010011001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10110010011001101011) && ({row_reg, col_reg}<20'b10110010100100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10110010100100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10110010100100011111) && ({row_reg, col_reg}<20'b10110010100101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10110010100101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10110010100101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10110010100101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10110010100101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10110010100101010000) && ({row_reg, col_reg}<20'b10110010101000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10110010101000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10110010101000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10110010101000111000) && ({row_reg, col_reg}<20'b10110010101000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10110010101000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10110010101000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10110010101000111100) && ({row_reg, col_reg}<20'b10110010101000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10110010101000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10110010101000111111) && ({row_reg, col_reg}<20'b10110010101001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10110010101001100110) && ({row_reg, col_reg}<20'b10110010101001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10110010101001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10110010101001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10110010101001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10110010101001101011) && ({row_reg, col_reg}<20'b10110010110100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10110010110100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10110010110100011111) && ({row_reg, col_reg}<20'b10110010110101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10110010110101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10110010110101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10110010110101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10110010110101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10110010110101010000) && ({row_reg, col_reg}<20'b10110010111000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10110010111000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10110010111000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10110010111000111000) && ({row_reg, col_reg}<20'b10110010111000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10110010111000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10110010111000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10110010111000111100) && ({row_reg, col_reg}<20'b10110010111000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10110010111000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10110010111000111111) && ({row_reg, col_reg}<20'b10110010111001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10110010111001100110) && ({row_reg, col_reg}<20'b10110010111001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10110010111001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10110010111001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10110010111001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10110010111001101011) && ({row_reg, col_reg}<20'b10110011000100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10110011000100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10110011000100011111) && ({row_reg, col_reg}<20'b10110011000101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10110011000101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10110011000101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10110011000101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10110011000101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10110011000101010000) && ({row_reg, col_reg}<20'b10110011001000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10110011001000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10110011001000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10110011001000111000) && ({row_reg, col_reg}<20'b10110011001000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10110011001000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10110011001000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10110011001000111100) && ({row_reg, col_reg}<20'b10110011001000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10110011001000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10110011001000111111) && ({row_reg, col_reg}<20'b10110011001001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10110011001001100110) && ({row_reg, col_reg}<20'b10110011001001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10110011001001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10110011001001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10110011001001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10110011001001101011) && ({row_reg, col_reg}<20'b10110011010100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10110011010100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10110011010100011111) && ({row_reg, col_reg}<20'b10110011010101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10110011010101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10110011010101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10110011010101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10110011010101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10110011010101010000) && ({row_reg, col_reg}<20'b10110011011000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10110011011000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10110011011000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10110011011000111000) && ({row_reg, col_reg}<20'b10110011011000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10110011011000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10110011011000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10110011011000111100) && ({row_reg, col_reg}<20'b10110011011000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10110011011000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10110011011000111111) && ({row_reg, col_reg}<20'b10110011011001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10110011011001100110) && ({row_reg, col_reg}<20'b10110011011001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10110011011001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10110011011001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10110011011001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10110011011001101011) && ({row_reg, col_reg}<20'b10110011100100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10110011100100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10110011100100011111) && ({row_reg, col_reg}<20'b10110011100101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10110011100101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10110011100101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10110011100101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10110011100101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10110011100101010000) && ({row_reg, col_reg}<20'b10110011101000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10110011101000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10110011101000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10110011101000111000) && ({row_reg, col_reg}<20'b10110011101000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10110011101000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10110011101000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10110011101000111100) && ({row_reg, col_reg}<20'b10110011101000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10110011101000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10110011101000111111) && ({row_reg, col_reg}<20'b10110011101001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10110011101001100110) && ({row_reg, col_reg}<20'b10110011101001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10110011101001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10110011101001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10110011101001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10110011101001101011) && ({row_reg, col_reg}<20'b10110011110100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10110011110100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10110011110100011111) && ({row_reg, col_reg}<20'b10110011110101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10110011110101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10110011110101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10110011110101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10110011110101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10110011110101010000) && ({row_reg, col_reg}<20'b10110011111000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10110011111000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10110011111000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10110011111000111000) && ({row_reg, col_reg}<20'b10110011111000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10110011111000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10110011111000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10110011111000111100) && ({row_reg, col_reg}<20'b10110011111000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10110011111000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10110011111000111111) && ({row_reg, col_reg}<20'b10110011111001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10110011111001100110) && ({row_reg, col_reg}<20'b10110011111001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10110011111001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10110011111001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10110011111001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10110011111001101011) && ({row_reg, col_reg}<20'b10110100000100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10110100000100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10110100000100011111) && ({row_reg, col_reg}<20'b10110100000101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10110100000101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10110100000101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10110100000101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10110100000101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10110100000101010000) && ({row_reg, col_reg}<20'b10110100001000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10110100001000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10110100001000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10110100001000111000) && ({row_reg, col_reg}<20'b10110100001000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10110100001000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10110100001000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10110100001000111100) && ({row_reg, col_reg}<20'b10110100001000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10110100001000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10110100001000111111) && ({row_reg, col_reg}<20'b10110100001001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10110100001001100110) && ({row_reg, col_reg}<20'b10110100001001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10110100001001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10110100001001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10110100001001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10110100001001101011) && ({row_reg, col_reg}<20'b10110100010100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10110100010100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10110100010100011111) && ({row_reg, col_reg}<20'b10110100010101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10110100010101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10110100010101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10110100010101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10110100010101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10110100010101010000) && ({row_reg, col_reg}<20'b10110100011000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10110100011000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10110100011000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10110100011000111000) && ({row_reg, col_reg}<20'b10110100011000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10110100011000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10110100011000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10110100011000111100) && ({row_reg, col_reg}<20'b10110100011000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10110100011000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10110100011000111111) && ({row_reg, col_reg}<20'b10110100011001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10110100011001100110) && ({row_reg, col_reg}<20'b10110100011001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10110100011001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10110100011001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10110100011001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10110100011001101011) && ({row_reg, col_reg}<20'b10110100100100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10110100100100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10110100100100011111) && ({row_reg, col_reg}<20'b10110100100101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10110100100101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10110100100101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10110100100101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10110100100101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10110100100101010000) && ({row_reg, col_reg}<20'b10110100101000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10110100101000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10110100101000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10110100101000111000) && ({row_reg, col_reg}<20'b10110100101000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10110100101000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10110100101000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10110100101000111100) && ({row_reg, col_reg}<20'b10110100101000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10110100101000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10110100101000111111) && ({row_reg, col_reg}<20'b10110100101001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10110100101001100110) && ({row_reg, col_reg}<20'b10110100101001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10110100101001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10110100101001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10110100101001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10110100101001101011) && ({row_reg, col_reg}<20'b10110100110100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10110100110100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10110100110100011111) && ({row_reg, col_reg}<20'b10110100110101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10110100110101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10110100110101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10110100110101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10110100110101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10110100110101010000) && ({row_reg, col_reg}<20'b10110100111000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10110100111000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10110100111000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10110100111000111000) && ({row_reg, col_reg}<20'b10110100111000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10110100111000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10110100111000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10110100111000111100) && ({row_reg, col_reg}<20'b10110100111000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10110100111000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10110100111000111111) && ({row_reg, col_reg}<20'b10110100111001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10110100111001100110) && ({row_reg, col_reg}<20'b10110100111001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10110100111001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10110100111001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10110100111001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10110100111001101011) && ({row_reg, col_reg}<20'b10110101000100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10110101000100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10110101000100011111) && ({row_reg, col_reg}<20'b10110101000101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10110101000101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10110101000101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10110101000101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10110101000101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10110101000101010000) && ({row_reg, col_reg}<20'b10110101001000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10110101001000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10110101001000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10110101001000111000) && ({row_reg, col_reg}<20'b10110101001000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10110101001000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10110101001000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10110101001000111100) && ({row_reg, col_reg}<20'b10110101001000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10110101001000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10110101001000111111) && ({row_reg, col_reg}<20'b10110101001001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10110101001001100110) && ({row_reg, col_reg}<20'b10110101001001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10110101001001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10110101001001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10110101001001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10110101001001101011) && ({row_reg, col_reg}<20'b10110101010100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10110101010100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10110101010100011111) && ({row_reg, col_reg}<20'b10110101010101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10110101010101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10110101010101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10110101010101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10110101010101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10110101010101010000) && ({row_reg, col_reg}<20'b10110101011000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10110101011000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10110101011000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10110101011000111000) && ({row_reg, col_reg}<20'b10110101011000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10110101011000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10110101011000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10110101011000111100) && ({row_reg, col_reg}<20'b10110101011000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10110101011000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10110101011000111111) && ({row_reg, col_reg}<20'b10110101011001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10110101011001100110) && ({row_reg, col_reg}<20'b10110101011001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10110101011001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10110101011001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10110101011001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10110101011001101011) && ({row_reg, col_reg}<20'b10110101100100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10110101100100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10110101100100011111) && ({row_reg, col_reg}<20'b10110101100101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10110101100101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10110101100101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10110101100101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10110101100101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10110101100101010000) && ({row_reg, col_reg}<20'b10110101101000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10110101101000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10110101101000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10110101101000111000) && ({row_reg, col_reg}<20'b10110101101000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10110101101000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10110101101000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10110101101000111100) && ({row_reg, col_reg}<20'b10110101101000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10110101101000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10110101101000111111) && ({row_reg, col_reg}<20'b10110101101001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10110101101001100110) && ({row_reg, col_reg}<20'b10110101101001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10110101101001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10110101101001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10110101101001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10110101101001101011) && ({row_reg, col_reg}<20'b10110101110100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10110101110100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10110101110100011111) && ({row_reg, col_reg}<20'b10110101110101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10110101110101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10110101110101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10110101110101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10110101110101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10110101110101010000) && ({row_reg, col_reg}<20'b10110101111000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10110101111000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10110101111000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10110101111000111000) && ({row_reg, col_reg}<20'b10110101111000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10110101111000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10110101111000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10110101111000111100) && ({row_reg, col_reg}<20'b10110101111000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10110101111000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10110101111000111111) && ({row_reg, col_reg}<20'b10110101111001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10110101111001100110) && ({row_reg, col_reg}<20'b10110101111001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10110101111001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10110101111001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10110101111001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10110101111001101011) && ({row_reg, col_reg}<20'b10110110000100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10110110000100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10110110000100011111) && ({row_reg, col_reg}<20'b10110110000101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10110110000101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10110110000101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10110110000101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10110110000101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10110110000101010000) && ({row_reg, col_reg}<20'b10110110001000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10110110001000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10110110001000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10110110001000111000) && ({row_reg, col_reg}<20'b10110110001000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10110110001000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10110110001000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10110110001000111100) && ({row_reg, col_reg}<20'b10110110001000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10110110001000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10110110001000111111) && ({row_reg, col_reg}<20'b10110110001001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10110110001001100110) && ({row_reg, col_reg}<20'b10110110001001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10110110001001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10110110001001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10110110001001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10110110001001101011) && ({row_reg, col_reg}<20'b10110110010100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10110110010100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10110110010100011111) && ({row_reg, col_reg}<20'b10110110010101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10110110010101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10110110010101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10110110010101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10110110010101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10110110010101010000) && ({row_reg, col_reg}<20'b10110110011000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10110110011000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10110110011000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10110110011000111000) && ({row_reg, col_reg}<20'b10110110011000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10110110011000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10110110011000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10110110011000111100) && ({row_reg, col_reg}<20'b10110110011000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10110110011000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10110110011000111111) && ({row_reg, col_reg}<20'b10110110011001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10110110011001100110) && ({row_reg, col_reg}<20'b10110110011001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10110110011001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10110110011001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10110110011001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10110110011001101011) && ({row_reg, col_reg}<20'b10110110100100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10110110100100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10110110100100011111) && ({row_reg, col_reg}<20'b10110110100101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10110110100101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10110110100101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10110110100101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10110110100101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10110110100101010000) && ({row_reg, col_reg}<20'b10110110101000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10110110101000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10110110101000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10110110101000111000) && ({row_reg, col_reg}<20'b10110110101000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10110110101000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10110110101000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10110110101000111100) && ({row_reg, col_reg}<20'b10110110101000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10110110101000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10110110101000111111) && ({row_reg, col_reg}<20'b10110110101001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10110110101001100110) && ({row_reg, col_reg}<20'b10110110101001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10110110101001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10110110101001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10110110101001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10110110101001101011) && ({row_reg, col_reg}<20'b10110110110100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10110110110100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10110110110100011111) && ({row_reg, col_reg}<20'b10110110110101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10110110110101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10110110110101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10110110110101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10110110110101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10110110110101010000) && ({row_reg, col_reg}<20'b10110110111000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10110110111000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10110110111000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10110110111000111000) && ({row_reg, col_reg}<20'b10110110111000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10110110111000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10110110111000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10110110111000111100) && ({row_reg, col_reg}<20'b10110110111000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10110110111000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10110110111000111111) && ({row_reg, col_reg}<20'b10110110111001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10110110111001100110) && ({row_reg, col_reg}<20'b10110110111001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10110110111001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10110110111001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10110110111001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10110110111001101011) && ({row_reg, col_reg}<20'b10110111000100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10110111000100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10110111000100011111) && ({row_reg, col_reg}<20'b10110111000101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10110111000101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10110111000101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10110111000101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10110111000101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10110111000101010000) && ({row_reg, col_reg}<20'b10110111001000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10110111001000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10110111001000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10110111001000111000) && ({row_reg, col_reg}<20'b10110111001000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10110111001000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10110111001000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10110111001000111100) && ({row_reg, col_reg}<20'b10110111001000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10110111001000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10110111001000111111) && ({row_reg, col_reg}<20'b10110111001001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10110111001001100110) && ({row_reg, col_reg}<20'b10110111001001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10110111001001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10110111001001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10110111001001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10110111001001101011) && ({row_reg, col_reg}<20'b10110111010100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10110111010100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10110111010100011111) && ({row_reg, col_reg}<20'b10110111010101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10110111010101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10110111010101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10110111010101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10110111010101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10110111010101010000) && ({row_reg, col_reg}<20'b10110111011000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10110111011000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10110111011000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10110111011000111000) && ({row_reg, col_reg}<20'b10110111011000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10110111011000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10110111011000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10110111011000111100) && ({row_reg, col_reg}<20'b10110111011000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10110111011000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10110111011000111111) && ({row_reg, col_reg}<20'b10110111011001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10110111011001100110) && ({row_reg, col_reg}<20'b10110111011001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10110111011001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10110111011001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10110111011001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10110111011001101011) && ({row_reg, col_reg}<20'b10110111100100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10110111100100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10110111100100011111) && ({row_reg, col_reg}<20'b10110111100101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10110111100101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10110111100101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10110111100101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10110111100101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10110111100101010000) && ({row_reg, col_reg}<20'b10110111101000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10110111101000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10110111101000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10110111101000111000) && ({row_reg, col_reg}<20'b10110111101000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10110111101000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10110111101000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10110111101000111100) && ({row_reg, col_reg}<20'b10110111101000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10110111101000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10110111101000111111) && ({row_reg, col_reg}<20'b10110111101001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10110111101001100110) && ({row_reg, col_reg}<20'b10110111101001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10110111101001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10110111101001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10110111101001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10110111101001101011) && ({row_reg, col_reg}<20'b10110111110100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10110111110100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10110111110100011111) && ({row_reg, col_reg}<20'b10110111110101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10110111110101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10110111110101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10110111110101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10110111110101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10110111110101010000) && ({row_reg, col_reg}<20'b10110111111000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10110111111000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10110111111000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10110111111000111000) && ({row_reg, col_reg}<20'b10110111111000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10110111111000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10110111111000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10110111111000111100) && ({row_reg, col_reg}<20'b10110111111000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10110111111000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10110111111000111111) && ({row_reg, col_reg}<20'b10110111111001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10110111111001100110) && ({row_reg, col_reg}<20'b10110111111001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10110111111001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10110111111001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10110111111001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10110111111001101011) && ({row_reg, col_reg}<20'b10111000000100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10111000000100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10111000000100011111) && ({row_reg, col_reg}<20'b10111000000101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10111000000101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10111000000101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10111000000101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10111000000101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10111000000101010000) && ({row_reg, col_reg}<20'b10111000001000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10111000001000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10111000001000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10111000001000111000) && ({row_reg, col_reg}<20'b10111000001000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10111000001000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10111000001000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10111000001000111100) && ({row_reg, col_reg}<20'b10111000001000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10111000001000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10111000001000111111) && ({row_reg, col_reg}<20'b10111000001001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10111000001001100110) && ({row_reg, col_reg}<20'b10111000001001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10111000001001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10111000001001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10111000001001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10111000001001101011) && ({row_reg, col_reg}<20'b10111000010100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10111000010100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10111000010100011111) && ({row_reg, col_reg}<20'b10111000010101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10111000010101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10111000010101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10111000010101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10111000010101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10111000010101010000) && ({row_reg, col_reg}<20'b10111000011000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10111000011000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10111000011000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10111000011000111000) && ({row_reg, col_reg}<20'b10111000011000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10111000011000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10111000011000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10111000011000111100) && ({row_reg, col_reg}<20'b10111000011000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10111000011000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10111000011000111111) && ({row_reg, col_reg}<20'b10111000011001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10111000011001100110) && ({row_reg, col_reg}<20'b10111000011001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10111000011001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10111000011001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10111000011001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10111000011001101011) && ({row_reg, col_reg}<20'b10111000100100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10111000100100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10111000100100011111) && ({row_reg, col_reg}<20'b10111000100101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10111000100101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10111000100101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10111000100101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10111000100101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10111000100101010000) && ({row_reg, col_reg}<20'b10111000101000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10111000101000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10111000101000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10111000101000111000) && ({row_reg, col_reg}<20'b10111000101000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10111000101000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10111000101000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10111000101000111100) && ({row_reg, col_reg}<20'b10111000101000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10111000101000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10111000101000111111) && ({row_reg, col_reg}<20'b10111000101001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10111000101001100110) && ({row_reg, col_reg}<20'b10111000101001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10111000101001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10111000101001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10111000101001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10111000101001101011) && ({row_reg, col_reg}<20'b10111000110100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10111000110100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10111000110100011111) && ({row_reg, col_reg}<20'b10111000110101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10111000110101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10111000110101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10111000110101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10111000110101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10111000110101010000) && ({row_reg, col_reg}<20'b10111000111000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10111000111000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10111000111000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10111000111000111000) && ({row_reg, col_reg}<20'b10111000111000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10111000111000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10111000111000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10111000111000111100) && ({row_reg, col_reg}<20'b10111000111000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10111000111000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10111000111000111111) && ({row_reg, col_reg}<20'b10111000111001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10111000111001100110) && ({row_reg, col_reg}<20'b10111000111001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10111000111001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10111000111001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10111000111001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10111000111001101011) && ({row_reg, col_reg}<20'b10111001000100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10111001000100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10111001000100011111) && ({row_reg, col_reg}<20'b10111001000101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10111001000101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10111001000101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10111001000101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10111001000101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10111001000101010000) && ({row_reg, col_reg}<20'b10111001001000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10111001001000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10111001001000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10111001001000111000) && ({row_reg, col_reg}<20'b10111001001000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10111001001000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10111001001000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10111001001000111100) && ({row_reg, col_reg}<20'b10111001001000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10111001001000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10111001001000111111) && ({row_reg, col_reg}<20'b10111001001001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10111001001001100110) && ({row_reg, col_reg}<20'b10111001001001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10111001001001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10111001001001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10111001001001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10111001001001101011) && ({row_reg, col_reg}<20'b10111001010100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10111001010100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10111001010100011111) && ({row_reg, col_reg}<20'b10111001010101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10111001010101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10111001010101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10111001010101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10111001010101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10111001010101010000) && ({row_reg, col_reg}<20'b10111001011000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10111001011000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10111001011000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10111001011000111000) && ({row_reg, col_reg}<20'b10111001011000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10111001011000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10111001011000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10111001011000111100) && ({row_reg, col_reg}<20'b10111001011000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10111001011000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10111001011000111111) && ({row_reg, col_reg}<20'b10111001011001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10111001011001100110) && ({row_reg, col_reg}<20'b10111001011001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10111001011001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10111001011001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10111001011001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10111001011001101011) && ({row_reg, col_reg}<20'b10111001100100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10111001100100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10111001100100011111) && ({row_reg, col_reg}<20'b10111001100101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10111001100101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10111001100101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10111001100101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10111001100101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10111001100101010000) && ({row_reg, col_reg}<20'b10111001101000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10111001101000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10111001101000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10111001101000111000) && ({row_reg, col_reg}<20'b10111001101000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10111001101000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10111001101000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10111001101000111100) && ({row_reg, col_reg}<20'b10111001101000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10111001101000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10111001101000111111) && ({row_reg, col_reg}<20'b10111001101001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10111001101001100110) && ({row_reg, col_reg}<20'b10111001101001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10111001101001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10111001101001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10111001101001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10111001101001101011) && ({row_reg, col_reg}<20'b10111001110100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10111001110100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10111001110100011111) && ({row_reg, col_reg}<20'b10111001110101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10111001110101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10111001110101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10111001110101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10111001110101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10111001110101010000) && ({row_reg, col_reg}<20'b10111001111000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10111001111000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10111001111000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10111001111000111000) && ({row_reg, col_reg}<20'b10111001111000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10111001111000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10111001111000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10111001111000111100) && ({row_reg, col_reg}<20'b10111001111000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10111001111000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10111001111000111111) && ({row_reg, col_reg}<20'b10111001111001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10111001111001100110) && ({row_reg, col_reg}<20'b10111001111001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10111001111001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10111001111001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10111001111001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10111001111001101011) && ({row_reg, col_reg}<20'b10111010000100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10111010000100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10111010000100011111) && ({row_reg, col_reg}<20'b10111010000101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10111010000101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10111010000101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10111010000101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10111010000101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10111010000101010000) && ({row_reg, col_reg}<20'b10111010001000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10111010001000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10111010001000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10111010001000111000) && ({row_reg, col_reg}<20'b10111010001000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10111010001000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10111010001000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10111010001000111100) && ({row_reg, col_reg}<20'b10111010001000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10111010001000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10111010001000111111) && ({row_reg, col_reg}<20'b10111010001001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10111010001001100110) && ({row_reg, col_reg}<20'b10111010001001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10111010001001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10111010001001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10111010001001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10111010001001101011) && ({row_reg, col_reg}<20'b10111010010100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10111010010100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10111010010100011111) && ({row_reg, col_reg}<20'b10111010010101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10111010010101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10111010010101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10111010010101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10111010010101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10111010010101010000) && ({row_reg, col_reg}<20'b10111010011000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10111010011000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10111010011000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10111010011000111000) && ({row_reg, col_reg}<20'b10111010011000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10111010011000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10111010011000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10111010011000111100) && ({row_reg, col_reg}<20'b10111010011000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10111010011000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10111010011000111111) && ({row_reg, col_reg}<20'b10111010011001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10111010011001100110) && ({row_reg, col_reg}<20'b10111010011001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10111010011001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10111010011001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10111010011001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10111010011001101011) && ({row_reg, col_reg}<20'b10111010100100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10111010100100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10111010100100011111) && ({row_reg, col_reg}<20'b10111010100101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10111010100101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10111010100101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10111010100101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10111010100101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10111010100101010000) && ({row_reg, col_reg}<20'b10111010101000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10111010101000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10111010101000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10111010101000111000) && ({row_reg, col_reg}<20'b10111010101000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10111010101000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10111010101000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10111010101000111100) && ({row_reg, col_reg}<20'b10111010101000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10111010101000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10111010101000111111) && ({row_reg, col_reg}<20'b10111010101001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10111010101001100110) && ({row_reg, col_reg}<20'b10111010101001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10111010101001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10111010101001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10111010101001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10111010101001101011) && ({row_reg, col_reg}<20'b10111010110100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10111010110100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10111010110100011111) && ({row_reg, col_reg}<20'b10111010110101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10111010110101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10111010110101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10111010110101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10111010110101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10111010110101010000) && ({row_reg, col_reg}<20'b10111010111000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10111010111000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10111010111000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10111010111000111000) && ({row_reg, col_reg}<20'b10111010111000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10111010111000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10111010111000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10111010111000111100) && ({row_reg, col_reg}<20'b10111010111000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10111010111000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10111010111000111111) && ({row_reg, col_reg}<20'b10111010111001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10111010111001100110) && ({row_reg, col_reg}<20'b10111010111001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10111010111001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10111010111001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10111010111001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10111010111001101011) && ({row_reg, col_reg}<20'b10111011000100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10111011000100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10111011000100011111) && ({row_reg, col_reg}<20'b10111011000101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10111011000101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10111011000101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10111011000101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10111011000101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10111011000101010000) && ({row_reg, col_reg}<20'b10111011001000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10111011001000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10111011001000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10111011001000111000) && ({row_reg, col_reg}<20'b10111011001000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10111011001000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10111011001000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10111011001000111100) && ({row_reg, col_reg}<20'b10111011001000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10111011001000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10111011001000111111) && ({row_reg, col_reg}<20'b10111011001001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10111011001001100110) && ({row_reg, col_reg}<20'b10111011001001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10111011001001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10111011001001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10111011001001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10111011001001101011) && ({row_reg, col_reg}<20'b10111011010100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10111011010100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10111011010100011111) && ({row_reg, col_reg}<20'b10111011010101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10111011010101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10111011010101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10111011010101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10111011010101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10111011010101010000) && ({row_reg, col_reg}<20'b10111011011000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10111011011000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10111011011000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10111011011000111000) && ({row_reg, col_reg}<20'b10111011011000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10111011011000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10111011011000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10111011011000111100) && ({row_reg, col_reg}<20'b10111011011000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10111011011000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10111011011000111111) && ({row_reg, col_reg}<20'b10111011011001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10111011011001100110) && ({row_reg, col_reg}<20'b10111011011001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10111011011001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10111011011001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10111011011001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10111011011001101011) && ({row_reg, col_reg}<20'b10111011100100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10111011100100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10111011100100011111) && ({row_reg, col_reg}<20'b10111011100101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10111011100101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10111011100101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10111011100101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10111011100101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10111011100101010000) && ({row_reg, col_reg}<20'b10111011101000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10111011101000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10111011101000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10111011101000111000) && ({row_reg, col_reg}<20'b10111011101000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10111011101000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10111011101000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10111011101000111100) && ({row_reg, col_reg}<20'b10111011101000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10111011101000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10111011101000111111) && ({row_reg, col_reg}<20'b10111011101001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10111011101001100110) && ({row_reg, col_reg}<20'b10111011101001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10111011101001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10111011101001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10111011101001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10111011101001101011) && ({row_reg, col_reg}<20'b10111011110100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10111011110100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10111011110100011111) && ({row_reg, col_reg}<20'b10111011110101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10111011110101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10111011110101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10111011110101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10111011110101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10111011110101010000) && ({row_reg, col_reg}<20'b10111011111000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10111011111000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10111011111000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10111011111000111000) && ({row_reg, col_reg}<20'b10111011111000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10111011111000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10111011111000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10111011111000111100) && ({row_reg, col_reg}<20'b10111011111000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10111011111000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10111011111000111111) && ({row_reg, col_reg}<20'b10111011111001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10111011111001100110) && ({row_reg, col_reg}<20'b10111011111001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10111011111001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10111011111001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10111011111001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10111011111001101011) && ({row_reg, col_reg}<20'b10111100000100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10111100000100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10111100000100011111) && ({row_reg, col_reg}<20'b10111100000101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10111100000101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10111100000101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10111100000101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10111100000101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10111100000101010000) && ({row_reg, col_reg}<20'b10111100001000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10111100001000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10111100001000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10111100001000111000) && ({row_reg, col_reg}<20'b10111100001000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10111100001000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10111100001000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10111100001000111100) && ({row_reg, col_reg}<20'b10111100001000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10111100001000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10111100001000111111) && ({row_reg, col_reg}<20'b10111100001001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10111100001001100110) && ({row_reg, col_reg}<20'b10111100001001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10111100001001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10111100001001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10111100001001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10111100001001101011) && ({row_reg, col_reg}<20'b10111100010100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10111100010100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10111100010100011111) && ({row_reg, col_reg}<20'b10111100010101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10111100010101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10111100010101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10111100010101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10111100010101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10111100010101010000) && ({row_reg, col_reg}<20'b10111100011000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10111100011000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10111100011000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10111100011000111000) && ({row_reg, col_reg}<20'b10111100011000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10111100011000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10111100011000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10111100011000111100) && ({row_reg, col_reg}<20'b10111100011000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10111100011000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10111100011000111111) && ({row_reg, col_reg}<20'b10111100011001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10111100011001100110) && ({row_reg, col_reg}<20'b10111100011001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10111100011001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10111100011001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10111100011001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10111100011001101011) && ({row_reg, col_reg}<20'b10111100100100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10111100100100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10111100100100011111) && ({row_reg, col_reg}<20'b10111100100101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10111100100101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10111100100101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10111100100101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10111100100101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10111100100101010000) && ({row_reg, col_reg}<20'b10111100101000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10111100101000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10111100101000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10111100101000111000) && ({row_reg, col_reg}<20'b10111100101000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10111100101000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10111100101000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10111100101000111100) && ({row_reg, col_reg}<20'b10111100101000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10111100101000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10111100101000111111) && ({row_reg, col_reg}<20'b10111100101001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10111100101001100110) && ({row_reg, col_reg}<20'b10111100101001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10111100101001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10111100101001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10111100101001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10111100101001101011) && ({row_reg, col_reg}<20'b10111100110100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10111100110100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10111100110100011111) && ({row_reg, col_reg}<20'b10111100110101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10111100110101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10111100110101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10111100110101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10111100110101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10111100110101010000) && ({row_reg, col_reg}<20'b10111100111000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10111100111000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10111100111000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10111100111000111000) && ({row_reg, col_reg}<20'b10111100111000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10111100111000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10111100111000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10111100111000111100) && ({row_reg, col_reg}<20'b10111100111000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10111100111000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10111100111000111111) && ({row_reg, col_reg}<20'b10111100111001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10111100111001100110) && ({row_reg, col_reg}<20'b10111100111001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10111100111001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10111100111001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10111100111001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10111100111001101011) && ({row_reg, col_reg}<20'b10111101000100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10111101000100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10111101000100011111) && ({row_reg, col_reg}<20'b10111101000101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10111101000101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10111101000101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10111101000101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10111101000101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10111101000101010000) && ({row_reg, col_reg}<20'b10111101001000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10111101001000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10111101001000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10111101001000111000) && ({row_reg, col_reg}<20'b10111101001000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10111101001000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10111101001000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10111101001000111100) && ({row_reg, col_reg}<20'b10111101001000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10111101001000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10111101001000111111) && ({row_reg, col_reg}<20'b10111101001001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10111101001001100110) && ({row_reg, col_reg}<20'b10111101001001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10111101001001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10111101001001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10111101001001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10111101001001101011) && ({row_reg, col_reg}<20'b10111101010100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10111101010100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10111101010100011111) && ({row_reg, col_reg}<20'b10111101010101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10111101010101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10111101010101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10111101010101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10111101010101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10111101010101010000) && ({row_reg, col_reg}<20'b10111101011000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10111101011000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10111101011000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10111101011000111000) && ({row_reg, col_reg}<20'b10111101011000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10111101011000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10111101011000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10111101011000111100) && ({row_reg, col_reg}<20'b10111101011000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10111101011000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10111101011000111111) && ({row_reg, col_reg}<20'b10111101011001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10111101011001100110) && ({row_reg, col_reg}<20'b10111101011001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10111101011001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10111101011001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10111101011001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10111101011001101011) && ({row_reg, col_reg}<20'b10111101100100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10111101100100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10111101100100011111) && ({row_reg, col_reg}<20'b10111101100101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10111101100101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10111101100101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10111101100101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10111101100101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10111101100101010000) && ({row_reg, col_reg}<20'b10111101101000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10111101101000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10111101101000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10111101101000111000) && ({row_reg, col_reg}<20'b10111101101000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10111101101000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10111101101000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10111101101000111100) && ({row_reg, col_reg}<20'b10111101101000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10111101101000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10111101101000111111) && ({row_reg, col_reg}<20'b10111101101001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10111101101001100110) && ({row_reg, col_reg}<20'b10111101101001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10111101101001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10111101101001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10111101101001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10111101101001101011) && ({row_reg, col_reg}<20'b10111101110100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10111101110100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10111101110100011111) && ({row_reg, col_reg}<20'b10111101110101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10111101110101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10111101110101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10111101110101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10111101110101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10111101110101010000) && ({row_reg, col_reg}<20'b10111101111000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10111101111000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10111101111000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10111101111000111000) && ({row_reg, col_reg}<20'b10111101111000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10111101111000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10111101111000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10111101111000111100) && ({row_reg, col_reg}<20'b10111101111000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10111101111000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10111101111000111111) && ({row_reg, col_reg}<20'b10111101111001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10111101111001100110) && ({row_reg, col_reg}<20'b10111101111001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10111101111001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10111101111001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10111101111001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10111101111001101011) && ({row_reg, col_reg}<20'b10111110000100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10111110000100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10111110000100011111) && ({row_reg, col_reg}<20'b10111110000101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10111110000101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10111110000101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10111110000101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10111110000101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10111110000101010000) && ({row_reg, col_reg}<20'b10111110001000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10111110001000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10111110001000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10111110001000111000) && ({row_reg, col_reg}<20'b10111110001000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10111110001000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10111110001000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10111110001000111100) && ({row_reg, col_reg}<20'b10111110001000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10111110001000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10111110001000111111) && ({row_reg, col_reg}<20'b10111110001001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10111110001001100110) && ({row_reg, col_reg}<20'b10111110001001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10111110001001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10111110001001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10111110001001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10111110001001101011) && ({row_reg, col_reg}<20'b10111110010100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10111110010100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10111110010100011111) && ({row_reg, col_reg}<20'b10111110010101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10111110010101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10111110010101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10111110010101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10111110010101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10111110010101010000) && ({row_reg, col_reg}<20'b10111110011000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10111110011000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10111110011000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10111110011000111000) && ({row_reg, col_reg}<20'b10111110011000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10111110011000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10111110011000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10111110011000111100) && ({row_reg, col_reg}<20'b10111110011000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10111110011000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10111110011000111111) && ({row_reg, col_reg}<20'b10111110011001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10111110011001100110) && ({row_reg, col_reg}<20'b10111110011001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10111110011001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10111110011001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10111110011001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10111110011001101011) && ({row_reg, col_reg}<20'b10111110100100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10111110100100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10111110100100011111) && ({row_reg, col_reg}<20'b10111110100101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10111110100101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10111110100101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10111110100101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10111110100101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10111110100101010000) && ({row_reg, col_reg}<20'b10111110101000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10111110101000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10111110101000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10111110101000111000) && ({row_reg, col_reg}<20'b10111110101000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10111110101000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10111110101000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10111110101000111100) && ({row_reg, col_reg}<20'b10111110101000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10111110101000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10111110101000111111) && ({row_reg, col_reg}<20'b10111110101001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10111110101001100110) && ({row_reg, col_reg}<20'b10111110101001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10111110101001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10111110101001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10111110101001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10111110101001101011) && ({row_reg, col_reg}<20'b10111110110100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10111110110100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10111110110100011111) && ({row_reg, col_reg}<20'b10111110110101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10111110110101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10111110110101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10111110110101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10111110110101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10111110110101010000) && ({row_reg, col_reg}<20'b10111110111000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10111110111000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10111110111000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10111110111000111000) && ({row_reg, col_reg}<20'b10111110111000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10111110111000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10111110111000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10111110111000111100) && ({row_reg, col_reg}<20'b10111110111000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10111110111000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10111110111000111111) && ({row_reg, col_reg}<20'b10111110111001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10111110111001100110) && ({row_reg, col_reg}<20'b10111110111001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10111110111001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10111110111001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10111110111001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10111110111001101011) && ({row_reg, col_reg}<20'b10111111000100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10111111000100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10111111000100011111) && ({row_reg, col_reg}<20'b10111111000101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10111111000101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10111111000101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10111111000101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10111111000101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10111111000101010000) && ({row_reg, col_reg}<20'b10111111001000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10111111001000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10111111001000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10111111001000111000) && ({row_reg, col_reg}<20'b10111111001000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10111111001000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10111111001000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10111111001000111100) && ({row_reg, col_reg}<20'b10111111001000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10111111001000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10111111001000111111) && ({row_reg, col_reg}<20'b10111111001001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10111111001001100110) && ({row_reg, col_reg}<20'b10111111001001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10111111001001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10111111001001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10111111001001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10111111001001101011) && ({row_reg, col_reg}<20'b10111111010100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10111111010100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10111111010100011111) && ({row_reg, col_reg}<20'b10111111010101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10111111010101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10111111010101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10111111010101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10111111010101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10111111010101010000) && ({row_reg, col_reg}<20'b10111111011000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10111111011000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10111111011000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10111111011000111000) && ({row_reg, col_reg}<20'b10111111011000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10111111011000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10111111011000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10111111011000111100) && ({row_reg, col_reg}<20'b10111111011000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10111111011000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10111111011000111111) && ({row_reg, col_reg}<20'b10111111011001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10111111011001100110) && ({row_reg, col_reg}<20'b10111111011001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10111111011001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10111111011001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10111111011001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10111111011001101011) && ({row_reg, col_reg}<20'b10111111100100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10111111100100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10111111100100011111) && ({row_reg, col_reg}<20'b10111111100101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10111111100101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10111111100101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10111111100101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10111111100101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10111111100101010000) && ({row_reg, col_reg}<20'b10111111101000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10111111101000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10111111101000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10111111101000111000) && ({row_reg, col_reg}<20'b10111111101000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10111111101000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10111111101000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10111111101000111100) && ({row_reg, col_reg}<20'b10111111101000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10111111101000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10111111101000111111) && ({row_reg, col_reg}<20'b10111111101001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10111111101001100110) && ({row_reg, col_reg}<20'b10111111101001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10111111101001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10111111101001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10111111101001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10111111101001101011) && ({row_reg, col_reg}<20'b10111111110100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10111111110100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b10111111110100011111) && ({row_reg, col_reg}<20'b10111111110101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10111111110101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10111111110101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10111111110101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10111111110101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10111111110101010000) && ({row_reg, col_reg}<20'b10111111111000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10111111111000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b10111111111000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b10111111111000111000) && ({row_reg, col_reg}<20'b10111111111000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10111111111000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10111111111000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10111111111000111100) && ({row_reg, col_reg}<20'b10111111111000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b10111111111000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b10111111111000111111) && ({row_reg, col_reg}<20'b10111111111001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b10111111111001100110) && ({row_reg, col_reg}<20'b10111111111001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b10111111111001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b10111111111001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b10111111111001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b10111111111001101011) && ({row_reg, col_reg}<20'b11000000000100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11000000000100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b11000000000100011111) && ({row_reg, col_reg}<20'b11000000000101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11000000000101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11000000000101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11000000000101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11000000000101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11000000000101010000) && ({row_reg, col_reg}<20'b11000000001000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11000000001000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b11000000001000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11000000001000111000) && ({row_reg, col_reg}<20'b11000000001000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11000000001000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11000000001000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11000000001000111100) && ({row_reg, col_reg}<20'b11000000001000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11000000001000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11000000001000111111) && ({row_reg, col_reg}<20'b11000000001001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b11000000001001100110) && ({row_reg, col_reg}<20'b11000000001001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11000000001001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b11000000001001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11000000001001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b11000000001001101011) && ({row_reg, col_reg}<20'b11000000010100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11000000010100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b11000000010100011111) && ({row_reg, col_reg}<20'b11000000010101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11000000010101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11000000010101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11000000010101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11000000010101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11000000010101010000) && ({row_reg, col_reg}<20'b11000000011000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11000000011000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b11000000011000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11000000011000111000) && ({row_reg, col_reg}<20'b11000000011000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11000000011000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11000000011000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11000000011000111100) && ({row_reg, col_reg}<20'b11000000011000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11000000011000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11000000011000111111) && ({row_reg, col_reg}<20'b11000000011001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b11000000011001100110) && ({row_reg, col_reg}<20'b11000000011001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11000000011001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b11000000011001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11000000011001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b11000000011001101011) && ({row_reg, col_reg}<20'b11000000100100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11000000100100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b11000000100100011111) && ({row_reg, col_reg}<20'b11000000100101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11000000100101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11000000100101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11000000100101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11000000100101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11000000100101010000) && ({row_reg, col_reg}<20'b11000000101000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11000000101000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b11000000101000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11000000101000111000) && ({row_reg, col_reg}<20'b11000000101000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11000000101000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11000000101000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11000000101000111100) && ({row_reg, col_reg}<20'b11000000101000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11000000101000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11000000101000111111) && ({row_reg, col_reg}<20'b11000000101001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b11000000101001100110) && ({row_reg, col_reg}<20'b11000000101001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11000000101001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b11000000101001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11000000101001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b11000000101001101011) && ({row_reg, col_reg}<20'b11000000110100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11000000110100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b11000000110100011111) && ({row_reg, col_reg}<20'b11000000110101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11000000110101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11000000110101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11000000110101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11000000110101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11000000110101010000) && ({row_reg, col_reg}<20'b11000000111000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11000000111000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b11000000111000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11000000111000111000) && ({row_reg, col_reg}<20'b11000000111000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11000000111000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11000000111000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11000000111000111100) && ({row_reg, col_reg}<20'b11000000111000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11000000111000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11000000111000111111) && ({row_reg, col_reg}<20'b11000000111001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b11000000111001100110) && ({row_reg, col_reg}<20'b11000000111001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11000000111001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b11000000111001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11000000111001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b11000000111001101011) && ({row_reg, col_reg}<20'b11000001000100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11000001000100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b11000001000100011111) && ({row_reg, col_reg}<20'b11000001000101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11000001000101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11000001000101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11000001000101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11000001000101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11000001000101010000) && ({row_reg, col_reg}<20'b11000001001000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11000001001000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b11000001001000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11000001001000111000) && ({row_reg, col_reg}<20'b11000001001000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11000001001000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11000001001000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11000001001000111100) && ({row_reg, col_reg}<20'b11000001001000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11000001001000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11000001001000111111) && ({row_reg, col_reg}<20'b11000001001001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b11000001001001100110) && ({row_reg, col_reg}<20'b11000001001001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11000001001001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b11000001001001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11000001001001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b11000001001001101011) && ({row_reg, col_reg}<20'b11000001010100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11000001010100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b11000001010100011111) && ({row_reg, col_reg}<20'b11000001010101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11000001010101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11000001010101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11000001010101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11000001010101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11000001010101010000) && ({row_reg, col_reg}<20'b11000001011000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11000001011000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b11000001011000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11000001011000111000) && ({row_reg, col_reg}<20'b11000001011000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11000001011000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11000001011000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11000001011000111100) && ({row_reg, col_reg}<20'b11000001011000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11000001011000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11000001011000111111) && ({row_reg, col_reg}<20'b11000001011001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b11000001011001100110) && ({row_reg, col_reg}<20'b11000001011001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11000001011001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b11000001011001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11000001011001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b11000001011001101011) && ({row_reg, col_reg}<20'b11000001100100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11000001100100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b11000001100100011111) && ({row_reg, col_reg}<20'b11000001100101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11000001100101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11000001100101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11000001100101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11000001100101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11000001100101010000) && ({row_reg, col_reg}<20'b11000001101000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11000001101000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b11000001101000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11000001101000111000) && ({row_reg, col_reg}<20'b11000001101000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11000001101000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11000001101000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11000001101000111100) && ({row_reg, col_reg}<20'b11000001101000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11000001101000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11000001101000111111) && ({row_reg, col_reg}<20'b11000001101001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b11000001101001100110) && ({row_reg, col_reg}<20'b11000001101001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11000001101001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b11000001101001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11000001101001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b11000001101001101011) && ({row_reg, col_reg}<20'b11000001110100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11000001110100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b11000001110100011111) && ({row_reg, col_reg}<20'b11000001110101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11000001110101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11000001110101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11000001110101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11000001110101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11000001110101010000) && ({row_reg, col_reg}<20'b11000001111000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11000001111000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b11000001111000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11000001111000111000) && ({row_reg, col_reg}<20'b11000001111000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11000001111000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11000001111000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11000001111000111100) && ({row_reg, col_reg}<20'b11000001111000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11000001111000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11000001111000111111) && ({row_reg, col_reg}<20'b11000001111001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b11000001111001100110) && ({row_reg, col_reg}<20'b11000001111001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11000001111001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b11000001111001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11000001111001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b11000001111001101011) && ({row_reg, col_reg}<20'b11000010000100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11000010000100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b11000010000100011111) && ({row_reg, col_reg}<20'b11000010000101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11000010000101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11000010000101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11000010000101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11000010000101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11000010000101010000) && ({row_reg, col_reg}<20'b11000010001000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11000010001000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b11000010001000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11000010001000111000) && ({row_reg, col_reg}<20'b11000010001000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11000010001000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11000010001000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11000010001000111100) && ({row_reg, col_reg}<20'b11000010001000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11000010001000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11000010001000111111) && ({row_reg, col_reg}<20'b11000010001001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b11000010001001100110) && ({row_reg, col_reg}<20'b11000010001001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11000010001001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b11000010001001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11000010001001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b11000010001001101011) && ({row_reg, col_reg}<20'b11000010010100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11000010010100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b11000010010100011111) && ({row_reg, col_reg}<20'b11000010010101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11000010010101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11000010010101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11000010010101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11000010010101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11000010010101010000) && ({row_reg, col_reg}<20'b11000010011000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11000010011000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b11000010011000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11000010011000111000) && ({row_reg, col_reg}<20'b11000010011000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11000010011000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11000010011000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11000010011000111100) && ({row_reg, col_reg}<20'b11000010011000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11000010011000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11000010011000111111) && ({row_reg, col_reg}<20'b11000010011001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b11000010011001100110) && ({row_reg, col_reg}<20'b11000010011001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11000010011001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b11000010011001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11000010011001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b11000010011001101011) && ({row_reg, col_reg}<20'b11000010100100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11000010100100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b11000010100100011111) && ({row_reg, col_reg}<20'b11000010100101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11000010100101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11000010100101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11000010100101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11000010100101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11000010100101010000) && ({row_reg, col_reg}<20'b11000010101000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11000010101000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b11000010101000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11000010101000111000) && ({row_reg, col_reg}<20'b11000010101000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11000010101000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11000010101000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11000010101000111100) && ({row_reg, col_reg}<20'b11000010101000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11000010101000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11000010101000111111) && ({row_reg, col_reg}<20'b11000010101001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b11000010101001100110) && ({row_reg, col_reg}<20'b11000010101001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11000010101001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b11000010101001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11000010101001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b11000010101001101011) && ({row_reg, col_reg}<20'b11000010110100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11000010110100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b11000010110100011111) && ({row_reg, col_reg}<20'b11000010110101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11000010110101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11000010110101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11000010110101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11000010110101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11000010110101010000) && ({row_reg, col_reg}<20'b11000010111000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11000010111000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b11000010111000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11000010111000111000) && ({row_reg, col_reg}<20'b11000010111000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11000010111000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11000010111000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11000010111000111100) && ({row_reg, col_reg}<20'b11000010111000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11000010111000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11000010111000111111) && ({row_reg, col_reg}<20'b11000010111001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b11000010111001100110) && ({row_reg, col_reg}<20'b11000010111001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11000010111001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b11000010111001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11000010111001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b11000010111001101011) && ({row_reg, col_reg}<20'b11000011000100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11000011000100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b11000011000100011111) && ({row_reg, col_reg}<20'b11000011000101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11000011000101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11000011000101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11000011000101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11000011000101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11000011000101010000) && ({row_reg, col_reg}<20'b11000011001000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11000011001000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b11000011001000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11000011001000111000) && ({row_reg, col_reg}<20'b11000011001000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11000011001000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11000011001000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11000011001000111100) && ({row_reg, col_reg}<20'b11000011001000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11000011001000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11000011001000111111) && ({row_reg, col_reg}<20'b11000011001001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b11000011001001100110) && ({row_reg, col_reg}<20'b11000011001001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11000011001001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b11000011001001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11000011001001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b11000011001001101011) && ({row_reg, col_reg}<20'b11000011010100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11000011010100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b11000011010100011111) && ({row_reg, col_reg}<20'b11000011010101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11000011010101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11000011010101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11000011010101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11000011010101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11000011010101010000) && ({row_reg, col_reg}<20'b11000011011000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11000011011000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b11000011011000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11000011011000111000) && ({row_reg, col_reg}<20'b11000011011000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11000011011000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11000011011000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11000011011000111100) && ({row_reg, col_reg}<20'b11000011011000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11000011011000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11000011011000111111) && ({row_reg, col_reg}<20'b11000011011001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b11000011011001100110) && ({row_reg, col_reg}<20'b11000011011001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11000011011001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b11000011011001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11000011011001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b11000011011001101011) && ({row_reg, col_reg}<20'b11000011100100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11000011100100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b11000011100100011111) && ({row_reg, col_reg}<20'b11000011100101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11000011100101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11000011100101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11000011100101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11000011100101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11000011100101010000) && ({row_reg, col_reg}<20'b11000011101000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11000011101000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b11000011101000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11000011101000111000) && ({row_reg, col_reg}<20'b11000011101000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11000011101000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11000011101000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11000011101000111100) && ({row_reg, col_reg}<20'b11000011101000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11000011101000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11000011101000111111) && ({row_reg, col_reg}<20'b11000011101001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b11000011101001100110) && ({row_reg, col_reg}<20'b11000011101001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11000011101001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b11000011101001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11000011101001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b11000011101001101011) && ({row_reg, col_reg}<20'b11000011110100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11000011110100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b11000011110100011111) && ({row_reg, col_reg}<20'b11000011110101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11000011110101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11000011110101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11000011110101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11000011110101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11000011110101010000) && ({row_reg, col_reg}<20'b11000011111000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11000011111000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b11000011111000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11000011111000111000) && ({row_reg, col_reg}<20'b11000011111000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11000011111000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11000011111000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11000011111000111100) && ({row_reg, col_reg}<20'b11000011111000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11000011111000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11000011111000111111) && ({row_reg, col_reg}<20'b11000011111001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b11000011111001100110) && ({row_reg, col_reg}<20'b11000011111001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11000011111001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b11000011111001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11000011111001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b11000011111001101011) && ({row_reg, col_reg}<20'b11000100000100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11000100000100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b11000100000100011111) && ({row_reg, col_reg}<20'b11000100000101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11000100000101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11000100000101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11000100000101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11000100000101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11000100000101010000) && ({row_reg, col_reg}<20'b11000100001000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11000100001000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b11000100001000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11000100001000111000) && ({row_reg, col_reg}<20'b11000100001000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11000100001000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11000100001000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11000100001000111100) && ({row_reg, col_reg}<20'b11000100001000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11000100001000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11000100001000111111) && ({row_reg, col_reg}<20'b11000100001001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b11000100001001100110) && ({row_reg, col_reg}<20'b11000100001001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11000100001001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b11000100001001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11000100001001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b11000100001001101011) && ({row_reg, col_reg}<20'b11000100010100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11000100010100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b11000100010100011111) && ({row_reg, col_reg}<20'b11000100010101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11000100010101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11000100010101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11000100010101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11000100010101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11000100010101010000) && ({row_reg, col_reg}<20'b11000100011000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11000100011000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b11000100011000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11000100011000111000) && ({row_reg, col_reg}<20'b11000100011000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11000100011000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11000100011000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11000100011000111100) && ({row_reg, col_reg}<20'b11000100011000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11000100011000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11000100011000111111) && ({row_reg, col_reg}<20'b11000100011001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b11000100011001100110) && ({row_reg, col_reg}<20'b11000100011001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11000100011001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b11000100011001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11000100011001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b11000100011001101011) && ({row_reg, col_reg}<20'b11000100100100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11000100100100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b11000100100100011111) && ({row_reg, col_reg}<20'b11000100100101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11000100100101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11000100100101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11000100100101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11000100100101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11000100100101010000) && ({row_reg, col_reg}<20'b11000100101000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11000100101000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b11000100101000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11000100101000111000) && ({row_reg, col_reg}<20'b11000100101000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11000100101000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11000100101000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11000100101000111100) && ({row_reg, col_reg}<20'b11000100101000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11000100101000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11000100101000111111) && ({row_reg, col_reg}<20'b11000100101001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b11000100101001100110) && ({row_reg, col_reg}<20'b11000100101001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11000100101001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b11000100101001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11000100101001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b11000100101001101011) && ({row_reg, col_reg}<20'b11000100110100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11000100110100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b11000100110100011111) && ({row_reg, col_reg}<20'b11000100110101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11000100110101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11000100110101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11000100110101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11000100110101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11000100110101010000) && ({row_reg, col_reg}<20'b11000100111000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11000100111000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b11000100111000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11000100111000111000) && ({row_reg, col_reg}<20'b11000100111000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11000100111000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11000100111000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11000100111000111100) && ({row_reg, col_reg}<20'b11000100111000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11000100111000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11000100111000111111) && ({row_reg, col_reg}<20'b11000100111001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b11000100111001100110) && ({row_reg, col_reg}<20'b11000100111001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11000100111001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b11000100111001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11000100111001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b11000100111001101011) && ({row_reg, col_reg}<20'b11000101000100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11000101000100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b11000101000100011111) && ({row_reg, col_reg}<20'b11000101000101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11000101000101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11000101000101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11000101000101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11000101000101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11000101000101010000) && ({row_reg, col_reg}<20'b11000101001000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11000101001000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b11000101001000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11000101001000111000) && ({row_reg, col_reg}<20'b11000101001000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11000101001000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11000101001000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11000101001000111100) && ({row_reg, col_reg}<20'b11000101001000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11000101001000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11000101001000111111) && ({row_reg, col_reg}<20'b11000101001001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b11000101001001100110) && ({row_reg, col_reg}<20'b11000101001001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11000101001001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b11000101001001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11000101001001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b11000101001001101011) && ({row_reg, col_reg}<20'b11000101010100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11000101010100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b11000101010100011111) && ({row_reg, col_reg}<20'b11000101010101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11000101010101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11000101010101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11000101010101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11000101010101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11000101010101010000) && ({row_reg, col_reg}<20'b11000101011000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11000101011000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b11000101011000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11000101011000111000) && ({row_reg, col_reg}<20'b11000101011000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11000101011000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11000101011000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11000101011000111100) && ({row_reg, col_reg}<20'b11000101011000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11000101011000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11000101011000111111) && ({row_reg, col_reg}<20'b11000101011001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b11000101011001100110) && ({row_reg, col_reg}<20'b11000101011001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11000101011001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b11000101011001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11000101011001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b11000101011001101011) && ({row_reg, col_reg}<20'b11000101100100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11000101100100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b11000101100100011111) && ({row_reg, col_reg}<20'b11000101100101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11000101100101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11000101100101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11000101100101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11000101100101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11000101100101010000) && ({row_reg, col_reg}<20'b11000101101000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11000101101000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b11000101101000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11000101101000111000) && ({row_reg, col_reg}<20'b11000101101000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11000101101000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11000101101000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11000101101000111100) && ({row_reg, col_reg}<20'b11000101101000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11000101101000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11000101101000111111) && ({row_reg, col_reg}<20'b11000101101001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b11000101101001100110) && ({row_reg, col_reg}<20'b11000101101001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11000101101001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b11000101101001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11000101101001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b11000101101001101011) && ({row_reg, col_reg}<20'b11000101110100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11000101110100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b11000101110100011111) && ({row_reg, col_reg}<20'b11000101110101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11000101110101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11000101110101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11000101110101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11000101110101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11000101110101010000) && ({row_reg, col_reg}<20'b11000101111000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11000101111000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b11000101111000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11000101111000111000) && ({row_reg, col_reg}<20'b11000101111000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11000101111000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11000101111000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11000101111000111100) && ({row_reg, col_reg}<20'b11000101111000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11000101111000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11000101111000111111) && ({row_reg, col_reg}<20'b11000101111001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b11000101111001100110) && ({row_reg, col_reg}<20'b11000101111001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11000101111001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b11000101111001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11000101111001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b11000101111001101011) && ({row_reg, col_reg}<20'b11000110000100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11000110000100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b11000110000100011111) && ({row_reg, col_reg}<20'b11000110000101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11000110000101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11000110000101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11000110000101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11000110000101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11000110000101010000) && ({row_reg, col_reg}<20'b11000110001000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11000110001000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b11000110001000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11000110001000111000) && ({row_reg, col_reg}<20'b11000110001000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11000110001000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11000110001000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11000110001000111100) && ({row_reg, col_reg}<20'b11000110001000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11000110001000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11000110001000111111) && ({row_reg, col_reg}<20'b11000110001001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b11000110001001100110) && ({row_reg, col_reg}<20'b11000110001001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11000110001001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b11000110001001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11000110001001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b11000110001001101011) && ({row_reg, col_reg}<20'b11000110010100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11000110010100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b11000110010100011111) && ({row_reg, col_reg}<20'b11000110010101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11000110010101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11000110010101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11000110010101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11000110010101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11000110010101010000) && ({row_reg, col_reg}<20'b11000110011000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11000110011000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b11000110011000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11000110011000111000) && ({row_reg, col_reg}<20'b11000110011000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11000110011000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11000110011000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11000110011000111100) && ({row_reg, col_reg}<20'b11000110011000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11000110011000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11000110011000111111) && ({row_reg, col_reg}<20'b11000110011001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b11000110011001100110) && ({row_reg, col_reg}<20'b11000110011001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11000110011001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b11000110011001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11000110011001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b11000110011001101011) && ({row_reg, col_reg}<20'b11000110100100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11000110100100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b11000110100100011111) && ({row_reg, col_reg}<20'b11000110100101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11000110100101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11000110100101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11000110100101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11000110100101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11000110100101010000) && ({row_reg, col_reg}<20'b11000110101000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11000110101000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b11000110101000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11000110101000111000) && ({row_reg, col_reg}<20'b11000110101000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11000110101000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11000110101000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11000110101000111100) && ({row_reg, col_reg}<20'b11000110101000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11000110101000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11000110101000111111) && ({row_reg, col_reg}<20'b11000110101001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b11000110101001100110) && ({row_reg, col_reg}<20'b11000110101001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11000110101001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b11000110101001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11000110101001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b11000110101001101011) && ({row_reg, col_reg}<20'b11000110110100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11000110110100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b11000110110100011111) && ({row_reg, col_reg}<20'b11000110110101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11000110110101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11000110110101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11000110110101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11000110110101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11000110110101010000) && ({row_reg, col_reg}<20'b11000110111000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11000110111000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b11000110111000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11000110111000111000) && ({row_reg, col_reg}<20'b11000110111000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11000110111000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11000110111000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11000110111000111100) && ({row_reg, col_reg}<20'b11000110111000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11000110111000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11000110111000111111) && ({row_reg, col_reg}<20'b11000110111001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b11000110111001100110) && ({row_reg, col_reg}<20'b11000110111001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11000110111001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b11000110111001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11000110111001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b11000110111001101011) && ({row_reg, col_reg}<20'b11000111000100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11000111000100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b11000111000100011111) && ({row_reg, col_reg}<20'b11000111000101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11000111000101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11000111000101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11000111000101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11000111000101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11000111000101010000) && ({row_reg, col_reg}<20'b11000111001000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11000111001000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b11000111001000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11000111001000111000) && ({row_reg, col_reg}<20'b11000111001000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11000111001000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11000111001000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11000111001000111100) && ({row_reg, col_reg}<20'b11000111001000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11000111001000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11000111001000111111) && ({row_reg, col_reg}<20'b11000111001001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b11000111001001100110) && ({row_reg, col_reg}<20'b11000111001001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11000111001001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b11000111001001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11000111001001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b11000111001001101011) && ({row_reg, col_reg}<20'b11000111010100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11000111010100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b11000111010100011111) && ({row_reg, col_reg}<20'b11000111010101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11000111010101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11000111010101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11000111010101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11000111010101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11000111010101010000) && ({row_reg, col_reg}<20'b11000111011000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11000111011000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b11000111011000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11000111011000111000) && ({row_reg, col_reg}<20'b11000111011000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11000111011000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11000111011000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11000111011000111100) && ({row_reg, col_reg}<20'b11000111011000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11000111011000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11000111011000111111) && ({row_reg, col_reg}<20'b11000111011001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b11000111011001100110) && ({row_reg, col_reg}<20'b11000111011001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11000111011001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b11000111011001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11000111011001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b11000111011001101011) && ({row_reg, col_reg}<20'b11000111100100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11000111100100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b11000111100100011111) && ({row_reg, col_reg}<20'b11000111100101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11000111100101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11000111100101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11000111100101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11000111100101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11000111100101010000) && ({row_reg, col_reg}<20'b11000111101000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11000111101000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b11000111101000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11000111101000111000) && ({row_reg, col_reg}<20'b11000111101000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11000111101000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11000111101000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11000111101000111100) && ({row_reg, col_reg}<20'b11000111101000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11000111101000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11000111101000111111) && ({row_reg, col_reg}<20'b11000111101001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b11000111101001100110) && ({row_reg, col_reg}<20'b11000111101001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11000111101001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b11000111101001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11000111101001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b11000111101001101011) && ({row_reg, col_reg}<20'b11000111110100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11000111110100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b11000111110100011111) && ({row_reg, col_reg}<20'b11000111110101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11000111110101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11000111110101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11000111110101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11000111110101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11000111110101010000) && ({row_reg, col_reg}<20'b11000111111000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11000111111000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b11000111111000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11000111111000111000) && ({row_reg, col_reg}<20'b11000111111000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11000111111000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11000111111000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11000111111000111100) && ({row_reg, col_reg}<20'b11000111111000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11000111111000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11000111111000111111) && ({row_reg, col_reg}<20'b11000111111001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b11000111111001100110) && ({row_reg, col_reg}<20'b11000111111001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11000111111001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b11000111111001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11000111111001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b11000111111001101011) && ({row_reg, col_reg}<20'b11001000000100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11001000000100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b11001000000100011111) && ({row_reg, col_reg}<20'b11001000000101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11001000000101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11001000000101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11001000000101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11001000000101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11001000000101010000) && ({row_reg, col_reg}<20'b11001000001000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11001000001000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b11001000001000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11001000001000111000) && ({row_reg, col_reg}<20'b11001000001000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11001000001000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11001000001000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11001000001000111100) && ({row_reg, col_reg}<20'b11001000001000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11001000001000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11001000001000111111) && ({row_reg, col_reg}<20'b11001000001001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b11001000001001100110) && ({row_reg, col_reg}<20'b11001000001001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11001000001001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b11001000001001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11001000001001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b11001000001001101011) && ({row_reg, col_reg}<20'b11001000010100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11001000010100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b11001000010100011111) && ({row_reg, col_reg}<20'b11001000010101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11001000010101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11001000010101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11001000010101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11001000010101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11001000010101010000) && ({row_reg, col_reg}<20'b11001000011000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11001000011000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b11001000011000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11001000011000111000) && ({row_reg, col_reg}<20'b11001000011000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11001000011000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11001000011000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11001000011000111100) && ({row_reg, col_reg}<20'b11001000011000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11001000011000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11001000011000111111) && ({row_reg, col_reg}<20'b11001000011001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b11001000011001100110) && ({row_reg, col_reg}<20'b11001000011001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11001000011001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b11001000011001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11001000011001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b11001000011001101011) && ({row_reg, col_reg}<20'b11001000100100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11001000100100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b11001000100100011111) && ({row_reg, col_reg}<20'b11001000100101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11001000100101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11001000100101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11001000100101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11001000100101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11001000100101010000) && ({row_reg, col_reg}<20'b11001000101000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11001000101000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b11001000101000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11001000101000111000) && ({row_reg, col_reg}<20'b11001000101000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11001000101000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11001000101000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11001000101000111100) && ({row_reg, col_reg}<20'b11001000101000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11001000101000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11001000101000111111) && ({row_reg, col_reg}<20'b11001000101001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b11001000101001100110) && ({row_reg, col_reg}<20'b11001000101001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11001000101001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b11001000101001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11001000101001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b11001000101001101011) && ({row_reg, col_reg}<20'b11001000110100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11001000110100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b11001000110100011111) && ({row_reg, col_reg}<20'b11001000110101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11001000110101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11001000110101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11001000110101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11001000110101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11001000110101010000) && ({row_reg, col_reg}<20'b11001000111000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11001000111000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b11001000111000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11001000111000111000) && ({row_reg, col_reg}<20'b11001000111000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11001000111000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11001000111000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11001000111000111100) && ({row_reg, col_reg}<20'b11001000111000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11001000111000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11001000111000111111) && ({row_reg, col_reg}<20'b11001000111001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b11001000111001100110) && ({row_reg, col_reg}<20'b11001000111001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11001000111001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b11001000111001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11001000111001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b11001000111001101011) && ({row_reg, col_reg}<20'b11001001000100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11001001000100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b11001001000100011111) && ({row_reg, col_reg}<20'b11001001000101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11001001000101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11001001000101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11001001000101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11001001000101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11001001000101010000) && ({row_reg, col_reg}<20'b11001001001000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11001001001000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b11001001001000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11001001001000111000) && ({row_reg, col_reg}<20'b11001001001000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11001001001000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11001001001000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11001001001000111100) && ({row_reg, col_reg}<20'b11001001001000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11001001001000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11001001001000111111) && ({row_reg, col_reg}<20'b11001001001001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b11001001001001100110) && ({row_reg, col_reg}<20'b11001001001001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11001001001001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b11001001001001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11001001001001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b11001001001001101011) && ({row_reg, col_reg}<20'b11001001010100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11001001010100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b11001001010100011111) && ({row_reg, col_reg}<20'b11001001010101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11001001010101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11001001010101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11001001010101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11001001010101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11001001010101010000) && ({row_reg, col_reg}<20'b11001001011000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11001001011000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b11001001011000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11001001011000111000) && ({row_reg, col_reg}<20'b11001001011000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11001001011000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11001001011000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11001001011000111100) && ({row_reg, col_reg}<20'b11001001011000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11001001011000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11001001011000111111) && ({row_reg, col_reg}<20'b11001001011001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b11001001011001100110) && ({row_reg, col_reg}<20'b11001001011001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11001001011001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b11001001011001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11001001011001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b11001001011001101011) && ({row_reg, col_reg}<20'b11001001100100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11001001100100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b11001001100100011111) && ({row_reg, col_reg}<20'b11001001100101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11001001100101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11001001100101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11001001100101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11001001100101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11001001100101010000) && ({row_reg, col_reg}<20'b11001001101000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11001001101000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b11001001101000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11001001101000111000) && ({row_reg, col_reg}<20'b11001001101000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11001001101000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11001001101000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11001001101000111100) && ({row_reg, col_reg}<20'b11001001101000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11001001101000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11001001101000111111) && ({row_reg, col_reg}<20'b11001001101001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b11001001101001100110) && ({row_reg, col_reg}<20'b11001001101001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11001001101001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b11001001101001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11001001101001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b11001001101001101011) && ({row_reg, col_reg}<20'b11001001110100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11001001110100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b11001001110100011111) && ({row_reg, col_reg}<20'b11001001110101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11001001110101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11001001110101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11001001110101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11001001110101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11001001110101010000) && ({row_reg, col_reg}<20'b11001001111000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11001001111000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b11001001111000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11001001111000111000) && ({row_reg, col_reg}<20'b11001001111000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11001001111000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11001001111000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11001001111000111100) && ({row_reg, col_reg}<20'b11001001111000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11001001111000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11001001111000111111) && ({row_reg, col_reg}<20'b11001001111001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b11001001111001100110) && ({row_reg, col_reg}<20'b11001001111001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11001001111001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b11001001111001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11001001111001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b11001001111001101011) && ({row_reg, col_reg}<20'b11001010000100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11001010000100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b11001010000100011111) && ({row_reg, col_reg}<20'b11001010000101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11001010000101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11001010000101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11001010000101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11001010000101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11001010000101010000) && ({row_reg, col_reg}<20'b11001010001000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11001010001000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b11001010001000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11001010001000111000) && ({row_reg, col_reg}<20'b11001010001000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11001010001000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11001010001000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11001010001000111100) && ({row_reg, col_reg}<20'b11001010001000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11001010001000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11001010001000111111) && ({row_reg, col_reg}<20'b11001010001001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b11001010001001100110) && ({row_reg, col_reg}<20'b11001010001001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11001010001001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b11001010001001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11001010001001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b11001010001001101011) && ({row_reg, col_reg}<20'b11001010010100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11001010010100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b11001010010100011111) && ({row_reg, col_reg}<20'b11001010010101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11001010010101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11001010010101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11001010010101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11001010010101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11001010010101010000) && ({row_reg, col_reg}<20'b11001010011000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11001010011000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b11001010011000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11001010011000111000) && ({row_reg, col_reg}<20'b11001010011000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11001010011000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11001010011000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11001010011000111100) && ({row_reg, col_reg}<20'b11001010011000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11001010011000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11001010011000111111) && ({row_reg, col_reg}<20'b11001010011001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b11001010011001100110) && ({row_reg, col_reg}<20'b11001010011001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11001010011001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b11001010011001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11001010011001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b11001010011001101011) && ({row_reg, col_reg}<20'b11001010100100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11001010100100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b11001010100100011111) && ({row_reg, col_reg}<20'b11001010100101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11001010100101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11001010100101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11001010100101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11001010100101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11001010100101010000) && ({row_reg, col_reg}<20'b11001010101000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11001010101000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b11001010101000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11001010101000111000) && ({row_reg, col_reg}<20'b11001010101000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11001010101000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11001010101000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11001010101000111100) && ({row_reg, col_reg}<20'b11001010101000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11001010101000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11001010101000111111) && ({row_reg, col_reg}<20'b11001010101001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b11001010101001100110) && ({row_reg, col_reg}<20'b11001010101001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11001010101001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b11001010101001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11001010101001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b11001010101001101011) && ({row_reg, col_reg}<20'b11001010110100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11001010110100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b11001010110100011111) && ({row_reg, col_reg}<20'b11001010110101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11001010110101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11001010110101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11001010110101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11001010110101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11001010110101010000) && ({row_reg, col_reg}<20'b11001010111000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11001010111000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b11001010111000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11001010111000111000) && ({row_reg, col_reg}<20'b11001010111000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11001010111000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11001010111000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11001010111000111100) && ({row_reg, col_reg}<20'b11001010111000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11001010111000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11001010111000111111) && ({row_reg, col_reg}<20'b11001010111001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b11001010111001100110) && ({row_reg, col_reg}<20'b11001010111001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11001010111001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b11001010111001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11001010111001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b11001010111001101011) && ({row_reg, col_reg}<20'b11001011000100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11001011000100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b11001011000100011111) && ({row_reg, col_reg}<20'b11001011000101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11001011000101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11001011000101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11001011000101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11001011000101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11001011000101010000) && ({row_reg, col_reg}<20'b11001011001000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11001011001000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b11001011001000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11001011001000111000) && ({row_reg, col_reg}<20'b11001011001000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11001011001000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11001011001000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11001011001000111100) && ({row_reg, col_reg}<20'b11001011001000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11001011001000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11001011001000111111) && ({row_reg, col_reg}<20'b11001011001001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b11001011001001100110) && ({row_reg, col_reg}<20'b11001011001001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11001011001001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b11001011001001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11001011001001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b11001011001001101011) && ({row_reg, col_reg}<20'b11001011010100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11001011010100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b11001011010100011111) && ({row_reg, col_reg}<20'b11001011010101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11001011010101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11001011010101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11001011010101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11001011010101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11001011010101010000) && ({row_reg, col_reg}<20'b11001011011000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11001011011000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b11001011011000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11001011011000111000) && ({row_reg, col_reg}<20'b11001011011000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11001011011000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11001011011000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11001011011000111100) && ({row_reg, col_reg}<20'b11001011011000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11001011011000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11001011011000111111) && ({row_reg, col_reg}<20'b11001011011001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b11001011011001100110) && ({row_reg, col_reg}<20'b11001011011001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11001011011001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b11001011011001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11001011011001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b11001011011001101011) && ({row_reg, col_reg}<20'b11001011100100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11001011100100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b11001011100100011111) && ({row_reg, col_reg}<20'b11001011100101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11001011100101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11001011100101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11001011100101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11001011100101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11001011100101010000) && ({row_reg, col_reg}<20'b11001011101000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11001011101000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b11001011101000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11001011101000111000) && ({row_reg, col_reg}<20'b11001011101000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11001011101000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11001011101000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11001011101000111100) && ({row_reg, col_reg}<20'b11001011101000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11001011101000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11001011101000111111) && ({row_reg, col_reg}<20'b11001011101001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b11001011101001100110) && ({row_reg, col_reg}<20'b11001011101001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11001011101001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b11001011101001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11001011101001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b11001011101001101011) && ({row_reg, col_reg}<20'b11001011110100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11001011110100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b11001011110100011111) && ({row_reg, col_reg}<20'b11001011110101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11001011110101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11001011110101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11001011110101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11001011110101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11001011110101010000) && ({row_reg, col_reg}<20'b11001011111000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11001011111000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b11001011111000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11001011111000111000) && ({row_reg, col_reg}<20'b11001011111000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11001011111000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11001011111000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11001011111000111100) && ({row_reg, col_reg}<20'b11001011111000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11001011111000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11001011111000111111) && ({row_reg, col_reg}<20'b11001011111001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b11001011111001100110) && ({row_reg, col_reg}<20'b11001011111001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11001011111001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b11001011111001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11001011111001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b11001011111001101011) && ({row_reg, col_reg}<20'b11001100000100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11001100000100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b11001100000100011111) && ({row_reg, col_reg}<20'b11001100000101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11001100000101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11001100000101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11001100000101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11001100000101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11001100000101010000) && ({row_reg, col_reg}<20'b11001100001000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11001100001000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b11001100001000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11001100001000111000) && ({row_reg, col_reg}<20'b11001100001000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11001100001000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11001100001000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11001100001000111100) && ({row_reg, col_reg}<20'b11001100001000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11001100001000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11001100001000111111) && ({row_reg, col_reg}<20'b11001100001001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b11001100001001100110) && ({row_reg, col_reg}<20'b11001100001001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11001100001001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b11001100001001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11001100001001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b11001100001001101011) && ({row_reg, col_reg}<20'b11001100010100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11001100010100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b11001100010100011111) && ({row_reg, col_reg}<20'b11001100010101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11001100010101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11001100010101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11001100010101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11001100010101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11001100010101010000) && ({row_reg, col_reg}<20'b11001100011000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11001100011000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b11001100011000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11001100011000111000) && ({row_reg, col_reg}<20'b11001100011000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11001100011000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11001100011000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11001100011000111100) && ({row_reg, col_reg}<20'b11001100011000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11001100011000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11001100011000111111) && ({row_reg, col_reg}<20'b11001100011001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b11001100011001100110) && ({row_reg, col_reg}<20'b11001100011001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11001100011001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b11001100011001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11001100011001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b11001100011001101011) && ({row_reg, col_reg}<20'b11001100100100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11001100100100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b11001100100100011111) && ({row_reg, col_reg}<20'b11001100100101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11001100100101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11001100100101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11001100100101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11001100100101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11001100100101010000) && ({row_reg, col_reg}<20'b11001100101000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11001100101000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b11001100101000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11001100101000111000) && ({row_reg, col_reg}<20'b11001100101000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11001100101000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11001100101000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11001100101000111100) && ({row_reg, col_reg}<20'b11001100101000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11001100101000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11001100101000111111) && ({row_reg, col_reg}<20'b11001100101001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b11001100101001100110) && ({row_reg, col_reg}<20'b11001100101001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11001100101001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b11001100101001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11001100101001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b11001100101001101011) && ({row_reg, col_reg}<20'b11001100110100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11001100110100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b11001100110100011111) && ({row_reg, col_reg}<20'b11001100110101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11001100110101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11001100110101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11001100110101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11001100110101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11001100110101010000) && ({row_reg, col_reg}<20'b11001100111000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11001100111000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b11001100111000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11001100111000111000) && ({row_reg, col_reg}<20'b11001100111000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11001100111000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11001100111000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11001100111000111100) && ({row_reg, col_reg}<20'b11001100111000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11001100111000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11001100111000111111) && ({row_reg, col_reg}<20'b11001100111001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b11001100111001100110) && ({row_reg, col_reg}<20'b11001100111001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11001100111001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b11001100111001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11001100111001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b11001100111001101011) && ({row_reg, col_reg}<20'b11001101000100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11001101000100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b11001101000100011111) && ({row_reg, col_reg}<20'b11001101000101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11001101000101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11001101000101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11001101000101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11001101000101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11001101000101010000) && ({row_reg, col_reg}<20'b11001101001000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11001101001000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b11001101001000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11001101001000111000) && ({row_reg, col_reg}<20'b11001101001000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11001101001000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11001101001000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11001101001000111100) && ({row_reg, col_reg}<20'b11001101001000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11001101001000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11001101001000111111) && ({row_reg, col_reg}<20'b11001101001001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b11001101001001100110) && ({row_reg, col_reg}<20'b11001101001001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11001101001001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b11001101001001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11001101001001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b11001101001001101011) && ({row_reg, col_reg}<20'b11001101010100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11001101010100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b11001101010100011111) && ({row_reg, col_reg}<20'b11001101010101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11001101010101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11001101010101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11001101010101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11001101010101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11001101010101010000) && ({row_reg, col_reg}<20'b11001101011000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11001101011000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b11001101011000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11001101011000111000) && ({row_reg, col_reg}<20'b11001101011000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11001101011000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11001101011000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11001101011000111100) && ({row_reg, col_reg}<20'b11001101011000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11001101011000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11001101011000111111) && ({row_reg, col_reg}<20'b11001101011001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b11001101011001100110) && ({row_reg, col_reg}<20'b11001101011001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11001101011001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b11001101011001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11001101011001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b11001101011001101011) && ({row_reg, col_reg}<20'b11001101100100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11001101100100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b11001101100100011111) && ({row_reg, col_reg}<20'b11001101100101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11001101100101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11001101100101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11001101100101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11001101100101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11001101100101010000) && ({row_reg, col_reg}<20'b11001101101000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11001101101000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b11001101101000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11001101101000111000) && ({row_reg, col_reg}<20'b11001101101000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11001101101000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11001101101000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11001101101000111100) && ({row_reg, col_reg}<20'b11001101101000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11001101101000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11001101101000111111) && ({row_reg, col_reg}<20'b11001101101001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b11001101101001100110) && ({row_reg, col_reg}<20'b11001101101001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11001101101001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b11001101101001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11001101101001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b11001101101001101011) && ({row_reg, col_reg}<20'b11001101110100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11001101110100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b11001101110100011111) && ({row_reg, col_reg}<20'b11001101110101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11001101110101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11001101110101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11001101110101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11001101110101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11001101110101010000) && ({row_reg, col_reg}<20'b11001101111000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11001101111000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b11001101111000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11001101111000111000) && ({row_reg, col_reg}<20'b11001101111000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11001101111000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11001101111000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11001101111000111100) && ({row_reg, col_reg}<20'b11001101111000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11001101111000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11001101111000111111) && ({row_reg, col_reg}<20'b11001101111001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b11001101111001100110) && ({row_reg, col_reg}<20'b11001101111001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11001101111001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b11001101111001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11001101111001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b11001101111001101011) && ({row_reg, col_reg}<20'b11001110000100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11001110000100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b11001110000100011111) && ({row_reg, col_reg}<20'b11001110000101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11001110000101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11001110000101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11001110000101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11001110000101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11001110000101010000) && ({row_reg, col_reg}<20'b11001110001000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11001110001000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b11001110001000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11001110001000111000) && ({row_reg, col_reg}<20'b11001110001000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11001110001000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11001110001000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11001110001000111100) && ({row_reg, col_reg}<20'b11001110001000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11001110001000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11001110001000111111) && ({row_reg, col_reg}<20'b11001110001001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b11001110001001100110) && ({row_reg, col_reg}<20'b11001110001001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11001110001001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b11001110001001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11001110001001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b11001110001001101011) && ({row_reg, col_reg}<20'b11001110010100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11001110010100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b11001110010100011111) && ({row_reg, col_reg}<20'b11001110010101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11001110010101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11001110010101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11001110010101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11001110010101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11001110010101010000) && ({row_reg, col_reg}<20'b11001110011000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11001110011000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b11001110011000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11001110011000111000) && ({row_reg, col_reg}<20'b11001110011000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11001110011000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11001110011000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11001110011000111100) && ({row_reg, col_reg}<20'b11001110011000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11001110011000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11001110011000111111) && ({row_reg, col_reg}<20'b11001110011001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b11001110011001100110) && ({row_reg, col_reg}<20'b11001110011001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11001110011001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b11001110011001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11001110011001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b11001110011001101011) && ({row_reg, col_reg}<20'b11001110100100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11001110100100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b11001110100100011111) && ({row_reg, col_reg}<20'b11001110100101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11001110100101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11001110100101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11001110100101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11001110100101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11001110100101010000) && ({row_reg, col_reg}<20'b11001110101000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11001110101000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b11001110101000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11001110101000111000) && ({row_reg, col_reg}<20'b11001110101000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11001110101000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11001110101000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11001110101000111100) && ({row_reg, col_reg}<20'b11001110101000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11001110101000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11001110101000111111) && ({row_reg, col_reg}<20'b11001110101001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b11001110101001100110) && ({row_reg, col_reg}<20'b11001110101001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11001110101001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b11001110101001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11001110101001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b11001110101001101011) && ({row_reg, col_reg}<20'b11001110110100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11001110110100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b11001110110100011111) && ({row_reg, col_reg}<20'b11001110110101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11001110110101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11001110110101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11001110110101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11001110110101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11001110110101010000) && ({row_reg, col_reg}<20'b11001110111000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11001110111000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b11001110111000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11001110111000111000) && ({row_reg, col_reg}<20'b11001110111000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11001110111000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11001110111000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11001110111000111100) && ({row_reg, col_reg}<20'b11001110111000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11001110111000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11001110111000111111) && ({row_reg, col_reg}<20'b11001110111001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b11001110111001100110) && ({row_reg, col_reg}<20'b11001110111001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11001110111001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b11001110111001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11001110111001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b11001110111001101011) && ({row_reg, col_reg}<20'b11001111000100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11001111000100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b11001111000100011111) && ({row_reg, col_reg}<20'b11001111000101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11001111000101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11001111000101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11001111000101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11001111000101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11001111000101010000) && ({row_reg, col_reg}<20'b11001111001000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11001111001000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b11001111001000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11001111001000111000) && ({row_reg, col_reg}<20'b11001111001000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11001111001000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11001111001000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11001111001000111100) && ({row_reg, col_reg}<20'b11001111001000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11001111001000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11001111001000111111) && ({row_reg, col_reg}<20'b11001111001001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b11001111001001100110) && ({row_reg, col_reg}<20'b11001111001001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11001111001001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b11001111001001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11001111001001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b11001111001001101011) && ({row_reg, col_reg}<20'b11001111010100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11001111010100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b11001111010100011111) && ({row_reg, col_reg}<20'b11001111010101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11001111010101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11001111010101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11001111010101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11001111010101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11001111010101010000) && ({row_reg, col_reg}<20'b11001111011000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11001111011000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b11001111011000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11001111011000111000) && ({row_reg, col_reg}<20'b11001111011000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11001111011000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11001111011000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11001111011000111100) && ({row_reg, col_reg}<20'b11001111011000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11001111011000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11001111011000111111) && ({row_reg, col_reg}<20'b11001111011001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b11001111011001100110) && ({row_reg, col_reg}<20'b11001111011001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11001111011001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b11001111011001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11001111011001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b11001111011001101011) && ({row_reg, col_reg}<20'b11001111100100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11001111100100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b11001111100100011111) && ({row_reg, col_reg}<20'b11001111100101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11001111100101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11001111100101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11001111100101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11001111100101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11001111100101010000) && ({row_reg, col_reg}<20'b11001111101000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11001111101000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b11001111101000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11001111101000111000) && ({row_reg, col_reg}<20'b11001111101000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11001111101000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11001111101000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11001111101000111100) && ({row_reg, col_reg}<20'b11001111101000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11001111101000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11001111101000111111) && ({row_reg, col_reg}<20'b11001111101001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b11001111101001100110) && ({row_reg, col_reg}<20'b11001111101001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11001111101001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b11001111101001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11001111101001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b11001111101001101011) && ({row_reg, col_reg}<20'b11001111110100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11001111110100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b11001111110100011111) && ({row_reg, col_reg}<20'b11001111110101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11001111110101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11001111110101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11001111110101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11001111110101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11001111110101010000) && ({row_reg, col_reg}<20'b11001111111000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11001111111000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b11001111111000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11001111111000111000) && ({row_reg, col_reg}<20'b11001111111000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11001111111000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11001111111000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11001111111000111100) && ({row_reg, col_reg}<20'b11001111111000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11001111111000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11001111111000111111) && ({row_reg, col_reg}<20'b11001111111001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b11001111111001100110) && ({row_reg, col_reg}<20'b11001111111001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11001111111001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b11001111111001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11001111111001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b11001111111001101011) && ({row_reg, col_reg}<20'b11010000000100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11010000000100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b11010000000100011111) && ({row_reg, col_reg}<20'b11010000000101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11010000000101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11010000000101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11010000000101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11010000000101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11010000000101010000) && ({row_reg, col_reg}<20'b11010000001000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11010000001000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b11010000001000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11010000001000111000) && ({row_reg, col_reg}<20'b11010000001000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11010000001000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11010000001000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11010000001000111100) && ({row_reg, col_reg}<20'b11010000001000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11010000001000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11010000001000111111) && ({row_reg, col_reg}<20'b11010000001001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b11010000001001100110) && ({row_reg, col_reg}<20'b11010000001001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11010000001001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b11010000001001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11010000001001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b11010000001001101011) && ({row_reg, col_reg}<20'b11010000010100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11010000010100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b11010000010100011111) && ({row_reg, col_reg}<20'b11010000010101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11010000010101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11010000010101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11010000010101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11010000010101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11010000010101010000) && ({row_reg, col_reg}<20'b11010000011000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11010000011000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b11010000011000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11010000011000111000) && ({row_reg, col_reg}<20'b11010000011000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11010000011000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11010000011000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11010000011000111100) && ({row_reg, col_reg}<20'b11010000011000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11010000011000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11010000011000111111) && ({row_reg, col_reg}<20'b11010000011001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b11010000011001100110) && ({row_reg, col_reg}<20'b11010000011001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11010000011001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b11010000011001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11010000011001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b11010000011001101011) && ({row_reg, col_reg}<20'b11010000100100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11010000100100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b11010000100100011111) && ({row_reg, col_reg}<20'b11010000100101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11010000100101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11010000100101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11010000100101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11010000100101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11010000100101010000) && ({row_reg, col_reg}<20'b11010000101000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11010000101000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b11010000101000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11010000101000111000) && ({row_reg, col_reg}<20'b11010000101000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11010000101000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11010000101000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11010000101000111100) && ({row_reg, col_reg}<20'b11010000101000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11010000101000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11010000101000111111) && ({row_reg, col_reg}<20'b11010000101001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b11010000101001100110) && ({row_reg, col_reg}<20'b11010000101001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11010000101001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b11010000101001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11010000101001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b11010000101001101011) && ({row_reg, col_reg}<20'b11010000110100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11010000110100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b11010000110100011111) && ({row_reg, col_reg}<20'b11010000110101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11010000110101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11010000110101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11010000110101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11010000110101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11010000110101010000) && ({row_reg, col_reg}<20'b11010000111000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11010000111000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b11010000111000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11010000111000111000) && ({row_reg, col_reg}<20'b11010000111000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11010000111000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11010000111000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11010000111000111100) && ({row_reg, col_reg}<20'b11010000111000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11010000111000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11010000111000111111) && ({row_reg, col_reg}<20'b11010000111001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b11010000111001100110) && ({row_reg, col_reg}<20'b11010000111001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11010000111001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b11010000111001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11010000111001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b11010000111001101011) && ({row_reg, col_reg}<20'b11010001000100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11010001000100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b11010001000100011111) && ({row_reg, col_reg}<20'b11010001000101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11010001000101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11010001000101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11010001000101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11010001000101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11010001000101010000) && ({row_reg, col_reg}<20'b11010001001000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11010001001000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b11010001001000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11010001001000111000) && ({row_reg, col_reg}<20'b11010001001000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11010001001000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11010001001000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11010001001000111100) && ({row_reg, col_reg}<20'b11010001001000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11010001001000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11010001001000111111) && ({row_reg, col_reg}<20'b11010001001001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b11010001001001100110) && ({row_reg, col_reg}<20'b11010001001001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11010001001001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b11010001001001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11010001001001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b11010001001001101011) && ({row_reg, col_reg}<20'b11010001010100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11010001010100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b11010001010100011111) && ({row_reg, col_reg}<20'b11010001010101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11010001010101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11010001010101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11010001010101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11010001010101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11010001010101010000) && ({row_reg, col_reg}<20'b11010001011000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11010001011000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b11010001011000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11010001011000111000) && ({row_reg, col_reg}<20'b11010001011000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11010001011000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11010001011000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11010001011000111100) && ({row_reg, col_reg}<20'b11010001011000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11010001011000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11010001011000111111) && ({row_reg, col_reg}<20'b11010001011001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b11010001011001100110) && ({row_reg, col_reg}<20'b11010001011001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11010001011001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b11010001011001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11010001011001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b11010001011001101011) && ({row_reg, col_reg}<20'b11010001100100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11010001100100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b11010001100100011111) && ({row_reg, col_reg}<20'b11010001100101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11010001100101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11010001100101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11010001100101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11010001100101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11010001100101010000) && ({row_reg, col_reg}<20'b11010001101000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11010001101000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b11010001101000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11010001101000111000) && ({row_reg, col_reg}<20'b11010001101000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11010001101000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11010001101000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11010001101000111100) && ({row_reg, col_reg}<20'b11010001101000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11010001101000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11010001101000111111) && ({row_reg, col_reg}<20'b11010001101001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b11010001101001100110) && ({row_reg, col_reg}<20'b11010001101001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11010001101001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b11010001101001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11010001101001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b11010001101001101011) && ({row_reg, col_reg}<20'b11010001110100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11010001110100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b11010001110100011111) && ({row_reg, col_reg}<20'b11010001110101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11010001110101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11010001110101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11010001110101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11010001110101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11010001110101010000) && ({row_reg, col_reg}<20'b11010001111000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11010001111000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b11010001111000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11010001111000111000) && ({row_reg, col_reg}<20'b11010001111000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11010001111000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11010001111000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11010001111000111100) && ({row_reg, col_reg}<20'b11010001111000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11010001111000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11010001111000111111) && ({row_reg, col_reg}<20'b11010001111001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b11010001111001100110) && ({row_reg, col_reg}<20'b11010001111001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11010001111001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b11010001111001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11010001111001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b11010001111001101011) && ({row_reg, col_reg}<20'b11010010000100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11010010000100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b11010010000100011111) && ({row_reg, col_reg}<20'b11010010000101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11010010000101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11010010000101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11010010000101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11010010000101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11010010000101010000) && ({row_reg, col_reg}<20'b11010010001000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11010010001000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b11010010001000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11010010001000111000) && ({row_reg, col_reg}<20'b11010010001000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11010010001000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11010010001000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11010010001000111100) && ({row_reg, col_reg}<20'b11010010001000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11010010001000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11010010001000111111) && ({row_reg, col_reg}<20'b11010010001001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b11010010001001100110) && ({row_reg, col_reg}<20'b11010010001001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11010010001001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b11010010001001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11010010001001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b11010010001001101011) && ({row_reg, col_reg}<20'b11010010010100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11010010010100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b11010010010100011111) && ({row_reg, col_reg}<20'b11010010010101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11010010010101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11010010010101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11010010010101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11010010010101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11010010010101010000) && ({row_reg, col_reg}<20'b11010010011000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11010010011000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b11010010011000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11010010011000111000) && ({row_reg, col_reg}<20'b11010010011000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11010010011000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11010010011000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11010010011000111100) && ({row_reg, col_reg}<20'b11010010011000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11010010011000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11010010011000111111) && ({row_reg, col_reg}<20'b11010010011001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b11010010011001100110) && ({row_reg, col_reg}<20'b11010010011001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11010010011001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b11010010011001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11010010011001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b11010010011001101011) && ({row_reg, col_reg}<20'b11010010100100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11010010100100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b11010010100100011111) && ({row_reg, col_reg}<20'b11010010100101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11010010100101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11010010100101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11010010100101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11010010100101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11010010100101010000) && ({row_reg, col_reg}<20'b11010010101000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11010010101000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b11010010101000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11010010101000111000) && ({row_reg, col_reg}<20'b11010010101000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11010010101000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11010010101000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11010010101000111100) && ({row_reg, col_reg}<20'b11010010101000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11010010101000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11010010101000111111) && ({row_reg, col_reg}<20'b11010010101001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b11010010101001100110) && ({row_reg, col_reg}<20'b11010010101001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11010010101001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b11010010101001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11010010101001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b11010010101001101011) && ({row_reg, col_reg}<20'b11010010110100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11010010110100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b11010010110100011111) && ({row_reg, col_reg}<20'b11010010110101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11010010110101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11010010110101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11010010110101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11010010110101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11010010110101010000) && ({row_reg, col_reg}<20'b11010010111000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11010010111000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b11010010111000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11010010111000111000) && ({row_reg, col_reg}<20'b11010010111000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11010010111000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11010010111000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11010010111000111100) && ({row_reg, col_reg}<20'b11010010111000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11010010111000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11010010111000111111) && ({row_reg, col_reg}<20'b11010010111001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b11010010111001100110) && ({row_reg, col_reg}<20'b11010010111001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11010010111001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b11010010111001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11010010111001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b11010010111001101011) && ({row_reg, col_reg}<20'b11010011000100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11010011000100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b11010011000100011111) && ({row_reg, col_reg}<20'b11010011000101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11010011000101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11010011000101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11010011000101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11010011000101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11010011000101010000) && ({row_reg, col_reg}<20'b11010011001000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11010011001000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b11010011001000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11010011001000111000) && ({row_reg, col_reg}<20'b11010011001000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11010011001000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11010011001000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11010011001000111100) && ({row_reg, col_reg}<20'b11010011001000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11010011001000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11010011001000111111) && ({row_reg, col_reg}<20'b11010011001001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b11010011001001100110) && ({row_reg, col_reg}<20'b11010011001001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11010011001001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b11010011001001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11010011001001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b11010011001001101011) && ({row_reg, col_reg}<20'b11010011010100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11010011010100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b11010011010100011111) && ({row_reg, col_reg}<20'b11010011010101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11010011010101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11010011010101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11010011010101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11010011010101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11010011010101010000) && ({row_reg, col_reg}<20'b11010011011000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11010011011000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b11010011011000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11010011011000111000) && ({row_reg, col_reg}<20'b11010011011000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11010011011000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11010011011000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11010011011000111100) && ({row_reg, col_reg}<20'b11010011011000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11010011011000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11010011011000111111) && ({row_reg, col_reg}<20'b11010011011001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b11010011011001100110) && ({row_reg, col_reg}<20'b11010011011001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11010011011001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b11010011011001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11010011011001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b11010011011001101011) && ({row_reg, col_reg}<20'b11010011100100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11010011100100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b11010011100100011111) && ({row_reg, col_reg}<20'b11010011100101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11010011100101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11010011100101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11010011100101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11010011100101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11010011100101010000) && ({row_reg, col_reg}<20'b11010011101000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11010011101000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b11010011101000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11010011101000111000) && ({row_reg, col_reg}<20'b11010011101000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11010011101000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11010011101000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11010011101000111100) && ({row_reg, col_reg}<20'b11010011101000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11010011101000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11010011101000111111) && ({row_reg, col_reg}<20'b11010011101001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b11010011101001100110) && ({row_reg, col_reg}<20'b11010011101001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11010011101001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b11010011101001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11010011101001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b11010011101001101011) && ({row_reg, col_reg}<20'b11010011110100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11010011110100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b11010011110100011111) && ({row_reg, col_reg}<20'b11010011110101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11010011110101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11010011110101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11010011110101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11010011110101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11010011110101010000) && ({row_reg, col_reg}<20'b11010011111000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11010011111000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b11010011111000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11010011111000111000) && ({row_reg, col_reg}<20'b11010011111000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11010011111000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11010011111000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11010011111000111100) && ({row_reg, col_reg}<20'b11010011111000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11010011111000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11010011111000111111) && ({row_reg, col_reg}<20'b11010011111001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b11010011111001100110) && ({row_reg, col_reg}<20'b11010011111001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11010011111001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b11010011111001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11010011111001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b11010011111001101011) && ({row_reg, col_reg}<20'b11010100000100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11010100000100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b11010100000100011111) && ({row_reg, col_reg}<20'b11010100000101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11010100000101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11010100000101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11010100000101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11010100000101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11010100000101010000) && ({row_reg, col_reg}<20'b11010100001000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11010100001000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b11010100001000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11010100001000111000) && ({row_reg, col_reg}<20'b11010100001000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11010100001000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11010100001000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11010100001000111100) && ({row_reg, col_reg}<20'b11010100001000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11010100001000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11010100001000111111) && ({row_reg, col_reg}<20'b11010100001001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b11010100001001100110) && ({row_reg, col_reg}<20'b11010100001001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11010100001001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b11010100001001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11010100001001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b11010100001001101011) && ({row_reg, col_reg}<20'b11010100010100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11010100010100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b11010100010100011111) && ({row_reg, col_reg}<20'b11010100010101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11010100010101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11010100010101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11010100010101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11010100010101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11010100010101010000) && ({row_reg, col_reg}<20'b11010100011000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11010100011000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b11010100011000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11010100011000111000) && ({row_reg, col_reg}<20'b11010100011000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11010100011000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11010100011000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11010100011000111100) && ({row_reg, col_reg}<20'b11010100011000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11010100011000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11010100011000111111) && ({row_reg, col_reg}<20'b11010100011001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b11010100011001100110) && ({row_reg, col_reg}<20'b11010100011001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11010100011001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b11010100011001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11010100011001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b11010100011001101011) && ({row_reg, col_reg}<20'b11010100100100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11010100100100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b11010100100100011111) && ({row_reg, col_reg}<20'b11010100100101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11010100100101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11010100100101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11010100100101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11010100100101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11010100100101010000) && ({row_reg, col_reg}<20'b11010100101000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11010100101000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b11010100101000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11010100101000111000) && ({row_reg, col_reg}<20'b11010100101000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11010100101000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11010100101000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11010100101000111100) && ({row_reg, col_reg}<20'b11010100101000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11010100101000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11010100101000111111) && ({row_reg, col_reg}<20'b11010100101001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b11010100101001100110) && ({row_reg, col_reg}<20'b11010100101001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11010100101001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b11010100101001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11010100101001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b11010100101001101011) && ({row_reg, col_reg}<20'b11010100110100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11010100110100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b11010100110100011111) && ({row_reg, col_reg}<20'b11010100110101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11010100110101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11010100110101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11010100110101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11010100110101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11010100110101010000) && ({row_reg, col_reg}<20'b11010100111000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11010100111000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b11010100111000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11010100111000111000) && ({row_reg, col_reg}<20'b11010100111000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11010100111000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11010100111000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11010100111000111100) && ({row_reg, col_reg}<20'b11010100111000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11010100111000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11010100111000111111) && ({row_reg, col_reg}<20'b11010100111001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b11010100111001100110) && ({row_reg, col_reg}<20'b11010100111001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11010100111001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b11010100111001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11010100111001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b11010100111001101011) && ({row_reg, col_reg}<20'b11010101000100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11010101000100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b11010101000100011111) && ({row_reg, col_reg}<20'b11010101000101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11010101000101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11010101000101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11010101000101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11010101000101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11010101000101010000) && ({row_reg, col_reg}<20'b11010101001000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11010101001000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b11010101001000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11010101001000111000) && ({row_reg, col_reg}<20'b11010101001000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11010101001000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11010101001000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11010101001000111100) && ({row_reg, col_reg}<20'b11010101001000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11010101001000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11010101001000111111) && ({row_reg, col_reg}<20'b11010101001001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b11010101001001100110) && ({row_reg, col_reg}<20'b11010101001001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11010101001001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b11010101001001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11010101001001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b11010101001001101011) && ({row_reg, col_reg}<20'b11010101010100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11010101010100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b11010101010100011111) && ({row_reg, col_reg}<20'b11010101010101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11010101010101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11010101010101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11010101010101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11010101010101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11010101010101010000) && ({row_reg, col_reg}<20'b11010101011000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11010101011000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b11010101011000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11010101011000111000) && ({row_reg, col_reg}<20'b11010101011000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11010101011000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11010101011000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11010101011000111100) && ({row_reg, col_reg}<20'b11010101011000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11010101011000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11010101011000111111) && ({row_reg, col_reg}<20'b11010101011001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b11010101011001100110) && ({row_reg, col_reg}<20'b11010101011001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11010101011001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b11010101011001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11010101011001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b11010101011001101011) && ({row_reg, col_reg}<20'b11010101100100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11010101100100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b11010101100100011111) && ({row_reg, col_reg}<20'b11010101100101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11010101100101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11010101100101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11010101100101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11010101100101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11010101100101010000) && ({row_reg, col_reg}<20'b11010101101000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11010101101000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b11010101101000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11010101101000111000) && ({row_reg, col_reg}<20'b11010101101000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11010101101000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11010101101000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11010101101000111100) && ({row_reg, col_reg}<20'b11010101101000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11010101101000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11010101101000111111) && ({row_reg, col_reg}<20'b11010101101001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b11010101101001100110) && ({row_reg, col_reg}<20'b11010101101001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11010101101001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b11010101101001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11010101101001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b11010101101001101011) && ({row_reg, col_reg}<20'b11010101110100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11010101110100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b11010101110100011111) && ({row_reg, col_reg}<20'b11010101110101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11010101110101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11010101110101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11010101110101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11010101110101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11010101110101010000) && ({row_reg, col_reg}<20'b11010101111000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11010101111000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b11010101111000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11010101111000111000) && ({row_reg, col_reg}<20'b11010101111000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11010101111000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11010101111000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11010101111000111100) && ({row_reg, col_reg}<20'b11010101111000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11010101111000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11010101111000111111) && ({row_reg, col_reg}<20'b11010101111001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b11010101111001100110) && ({row_reg, col_reg}<20'b11010101111001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11010101111001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b11010101111001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11010101111001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b11010101111001101011) && ({row_reg, col_reg}<20'b11010110000100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11010110000100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b11010110000100011111) && ({row_reg, col_reg}<20'b11010110000101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11010110000101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11010110000101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11010110000101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11010110000101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11010110000101010000) && ({row_reg, col_reg}<20'b11010110001000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11010110001000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b11010110001000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11010110001000111000) && ({row_reg, col_reg}<20'b11010110001000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11010110001000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11010110001000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11010110001000111100) && ({row_reg, col_reg}<20'b11010110001000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11010110001000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11010110001000111111) && ({row_reg, col_reg}<20'b11010110001001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b11010110001001100110) && ({row_reg, col_reg}<20'b11010110001001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11010110001001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b11010110001001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11010110001001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b11010110001001101011) && ({row_reg, col_reg}<20'b11010110010100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11010110010100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b11010110010100011111) && ({row_reg, col_reg}<20'b11010110010101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11010110010101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11010110010101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11010110010101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11010110010101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11010110010101010000) && ({row_reg, col_reg}<20'b11010110011000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11010110011000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b11010110011000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11010110011000111000) && ({row_reg, col_reg}<20'b11010110011000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11010110011000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11010110011000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11010110011000111100) && ({row_reg, col_reg}<20'b11010110011000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11010110011000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11010110011000111111) && ({row_reg, col_reg}<20'b11010110011001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b11010110011001100110) && ({row_reg, col_reg}<20'b11010110011001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11010110011001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b11010110011001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11010110011001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b11010110011001101011) && ({row_reg, col_reg}<20'b11010110100100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11010110100100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b11010110100100011111) && ({row_reg, col_reg}<20'b11010110100101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11010110100101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11010110100101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11010110100101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11010110100101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11010110100101010000) && ({row_reg, col_reg}<20'b11010110101000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11010110101000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b11010110101000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11010110101000111000) && ({row_reg, col_reg}<20'b11010110101000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11010110101000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11010110101000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11010110101000111100) && ({row_reg, col_reg}<20'b11010110101000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11010110101000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11010110101000111111) && ({row_reg, col_reg}<20'b11010110101001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b11010110101001100110) && ({row_reg, col_reg}<20'b11010110101001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11010110101001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b11010110101001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11010110101001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b11010110101001101011) && ({row_reg, col_reg}<20'b11010110110100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11010110110100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b11010110110100011111) && ({row_reg, col_reg}<20'b11010110110101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11010110110101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11010110110101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11010110110101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11010110110101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11010110110101010000) && ({row_reg, col_reg}<20'b11010110111000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11010110111000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b11010110111000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11010110111000111000) && ({row_reg, col_reg}<20'b11010110111000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11010110111000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11010110111000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11010110111000111100) && ({row_reg, col_reg}<20'b11010110111000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11010110111000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11010110111000111111) && ({row_reg, col_reg}<20'b11010110111001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b11010110111001100110) && ({row_reg, col_reg}<20'b11010110111001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11010110111001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b11010110111001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11010110111001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b11010110111001101011) && ({row_reg, col_reg}<20'b11010111000100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11010111000100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b11010111000100011111) && ({row_reg, col_reg}<20'b11010111000101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11010111000101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11010111000101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11010111000101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11010111000101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11010111000101010000) && ({row_reg, col_reg}<20'b11010111001000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11010111001000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b11010111001000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11010111001000111000) && ({row_reg, col_reg}<20'b11010111001000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11010111001000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11010111001000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11010111001000111100) && ({row_reg, col_reg}<20'b11010111001000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11010111001000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11010111001000111111) && ({row_reg, col_reg}<20'b11010111001001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b11010111001001100110) && ({row_reg, col_reg}<20'b11010111001001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11010111001001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b11010111001001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11010111001001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b11010111001001101011) && ({row_reg, col_reg}<20'b11010111010100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11010111010100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b11010111010100011111) && ({row_reg, col_reg}<20'b11010111010101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11010111010101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11010111010101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11010111010101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11010111010101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11010111010101010000) && ({row_reg, col_reg}<20'b11010111011000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11010111011000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b11010111011000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11010111011000111000) && ({row_reg, col_reg}<20'b11010111011000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11010111011000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11010111011000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11010111011000111100) && ({row_reg, col_reg}<20'b11010111011000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11010111011000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11010111011000111111) && ({row_reg, col_reg}<20'b11010111011001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b11010111011001100110) && ({row_reg, col_reg}<20'b11010111011001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11010111011001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b11010111011001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11010111011001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b11010111011001101011) && ({row_reg, col_reg}<20'b11010111100100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11010111100100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b11010111100100011111) && ({row_reg, col_reg}<20'b11010111100101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11010111100101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11010111100101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11010111100101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11010111100101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11010111100101010000) && ({row_reg, col_reg}<20'b11010111101000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11010111101000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b11010111101000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11010111101000111000) && ({row_reg, col_reg}<20'b11010111101000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11010111101000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11010111101000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11010111101000111100) && ({row_reg, col_reg}<20'b11010111101000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11010111101000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11010111101000111111) && ({row_reg, col_reg}<20'b11010111101001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b11010111101001100110) && ({row_reg, col_reg}<20'b11010111101001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11010111101001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b11010111101001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11010111101001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b11010111101001101011) && ({row_reg, col_reg}<20'b11010111110100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11010111110100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b11010111110100011111) && ({row_reg, col_reg}<20'b11010111110101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11010111110101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11010111110101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11010111110101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11010111110101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11010111110101010000) && ({row_reg, col_reg}<20'b11010111111000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11010111111000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b11010111111000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11010111111000111000) && ({row_reg, col_reg}<20'b11010111111000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11010111111000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11010111111000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11010111111000111100) && ({row_reg, col_reg}<20'b11010111111000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11010111111000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11010111111000111111) && ({row_reg, col_reg}<20'b11010111111001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b11010111111001100110) && ({row_reg, col_reg}<20'b11010111111001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11010111111001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b11010111111001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11010111111001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b11010111111001101011) && ({row_reg, col_reg}<20'b11011000000100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11011000000100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b11011000000100011111) && ({row_reg, col_reg}<20'b11011000000101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11011000000101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11011000000101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11011000000101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11011000000101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11011000000101010000) && ({row_reg, col_reg}<20'b11011000001000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11011000001000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b11011000001000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11011000001000111000) && ({row_reg, col_reg}<20'b11011000001000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11011000001000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11011000001000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11011000001000111100) && ({row_reg, col_reg}<20'b11011000001000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11011000001000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11011000001000111111) && ({row_reg, col_reg}<20'b11011000001001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b11011000001001100110) && ({row_reg, col_reg}<20'b11011000001001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11011000001001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b11011000001001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11011000001001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b11011000001001101011) && ({row_reg, col_reg}<20'b11011000010100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11011000010100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b11011000010100011111) && ({row_reg, col_reg}<20'b11011000010101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11011000010101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11011000010101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11011000010101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11011000010101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11011000010101010000) && ({row_reg, col_reg}<20'b11011000011000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11011000011000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b11011000011000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11011000011000111000) && ({row_reg, col_reg}<20'b11011000011000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11011000011000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11011000011000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11011000011000111100) && ({row_reg, col_reg}<20'b11011000011000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11011000011000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11011000011000111111) && ({row_reg, col_reg}<20'b11011000011001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b11011000011001100110) && ({row_reg, col_reg}<20'b11011000011001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11011000011001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b11011000011001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11011000011001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b11011000011001101011) && ({row_reg, col_reg}<20'b11011000100100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11011000100100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b11011000100100011111) && ({row_reg, col_reg}<20'b11011000100101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11011000100101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11011000100101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11011000100101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11011000100101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11011000100101010000) && ({row_reg, col_reg}<20'b11011000101000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11011000101000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b11011000101000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11011000101000111000) && ({row_reg, col_reg}<20'b11011000101000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11011000101000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11011000101000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11011000101000111100) && ({row_reg, col_reg}<20'b11011000101000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11011000101000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11011000101000111111) && ({row_reg, col_reg}<20'b11011000101001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b11011000101001100110) && ({row_reg, col_reg}<20'b11011000101001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11011000101001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b11011000101001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11011000101001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b11011000101001101011) && ({row_reg, col_reg}<20'b11011000110100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11011000110100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b11011000110100011111) && ({row_reg, col_reg}<20'b11011000110101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11011000110101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11011000110101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11011000110101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11011000110101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11011000110101010000) && ({row_reg, col_reg}<20'b11011000111000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11011000111000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b11011000111000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11011000111000111000) && ({row_reg, col_reg}<20'b11011000111000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11011000111000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11011000111000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11011000111000111100) && ({row_reg, col_reg}<20'b11011000111000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11011000111000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11011000111000111111) && ({row_reg, col_reg}<20'b11011000111001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b11011000111001100110) && ({row_reg, col_reg}<20'b11011000111001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11011000111001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b11011000111001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11011000111001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b11011000111001101011) && ({row_reg, col_reg}<20'b11011001000100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11011001000100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b11011001000100011111) && ({row_reg, col_reg}<20'b11011001000101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11011001000101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11011001000101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11011001000101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11011001000101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11011001000101010000) && ({row_reg, col_reg}<20'b11011001001000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11011001001000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b11011001001000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11011001001000111000) && ({row_reg, col_reg}<20'b11011001001000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11011001001000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11011001001000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11011001001000111100) && ({row_reg, col_reg}<20'b11011001001000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11011001001000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11011001001000111111) && ({row_reg, col_reg}<20'b11011001001001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b11011001001001100110) && ({row_reg, col_reg}<20'b11011001001001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11011001001001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b11011001001001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11011001001001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b11011001001001101011) && ({row_reg, col_reg}<20'b11011001010100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11011001010100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b11011001010100011111) && ({row_reg, col_reg}<20'b11011001010101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11011001010101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11011001010101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11011001010101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11011001010101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11011001010101010000) && ({row_reg, col_reg}<20'b11011001011000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11011001011000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b11011001011000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11011001011000111000) && ({row_reg, col_reg}<20'b11011001011000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11011001011000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11011001011000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11011001011000111100) && ({row_reg, col_reg}<20'b11011001011000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11011001011000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11011001011000111111) && ({row_reg, col_reg}<20'b11011001011001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b11011001011001100110) && ({row_reg, col_reg}<20'b11011001011001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11011001011001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b11011001011001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11011001011001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b11011001011001101011) && ({row_reg, col_reg}<20'b11011001100100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11011001100100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b11011001100100011111) && ({row_reg, col_reg}<20'b11011001100101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11011001100101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11011001100101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11011001100101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11011001100101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11011001100101010000) && ({row_reg, col_reg}<20'b11011001101000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11011001101000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b11011001101000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11011001101000111000) && ({row_reg, col_reg}<20'b11011001101000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11011001101000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11011001101000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11011001101000111100) && ({row_reg, col_reg}<20'b11011001101000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11011001101000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11011001101000111111) && ({row_reg, col_reg}<20'b11011001101001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b11011001101001100110) && ({row_reg, col_reg}<20'b11011001101001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11011001101001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b11011001101001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11011001101001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b11011001101001101011) && ({row_reg, col_reg}<20'b11011001110100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11011001110100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b11011001110100011111) && ({row_reg, col_reg}<20'b11011001110101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11011001110101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11011001110101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11011001110101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11011001110101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11011001110101010000) && ({row_reg, col_reg}<20'b11011001111000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11011001111000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b11011001111000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11011001111000111000) && ({row_reg, col_reg}<20'b11011001111000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11011001111000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11011001111000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11011001111000111100) && ({row_reg, col_reg}<20'b11011001111000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11011001111000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11011001111000111111) && ({row_reg, col_reg}<20'b11011001111001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b11011001111001100110) && ({row_reg, col_reg}<20'b11011001111001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11011001111001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b11011001111001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11011001111001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b11011001111001101011) && ({row_reg, col_reg}<20'b11011010000100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11011010000100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b11011010000100011111) && ({row_reg, col_reg}<20'b11011010000101001001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11011010000101001001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11011010000101001010) && ({row_reg, col_reg}<20'b11011010000101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11011010000101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11011010000101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11011010000101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11011010000101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11011010000101010000) && ({row_reg, col_reg}<20'b11011010001000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11011010001000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b11011010001000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11011010001000111000) && ({row_reg, col_reg}<20'b11011010001000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11011010001000111010) && ({row_reg, col_reg}<20'b11011010001000111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11011010001000111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11011010001000111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11011010001000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11011010001000111111) && ({row_reg, col_reg}<20'b11011010001001100000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11011010001001100000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11011010001001100001) && ({row_reg, col_reg}<20'b11011010001001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b11011010001001100110) && ({row_reg, col_reg}<20'b11011010001001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11011010001001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b11011010001001101001) && ({row_reg, col_reg}<20'b11011010001001101100)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11011010001001101100)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b11011010001001101101) && ({row_reg, col_reg}<20'b11011010010100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11011010010100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b11011010010100011111) && ({row_reg, col_reg}<20'b11011010010101001001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11011010010101001001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11011010010101001010) && ({row_reg, col_reg}<20'b11011010010101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11011010010101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11011010010101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11011010010101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11011010010101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11011010010101010000) && ({row_reg, col_reg}<20'b11011010011000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11011010011000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b11011010011000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11011010011000111000) && ({row_reg, col_reg}<20'b11011010011000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11011010011000111010) && ({row_reg, col_reg}<20'b11011010011000111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11011010011000111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11011010011000111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11011010011000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11011010011000111111) && ({row_reg, col_reg}<20'b11011010011001100000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11011010011001100000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11011010011001100001) && ({row_reg, col_reg}<20'b11011010011001100101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b11011010011001100101) && ({row_reg, col_reg}<20'b11011010011001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11011010011001101000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b11011010011001101001) && ({row_reg, col_reg}<20'b11011010011001101100)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11011010011001101100)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b11011010011001101101) && ({row_reg, col_reg}<20'b11011010100100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11011010100100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b11011010100100011111) && ({row_reg, col_reg}<20'b11011010100101001001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11011010100101001001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11011010100101001010) && ({row_reg, col_reg}<20'b11011010100101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11011010100101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11011010100101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11011010100101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11011010100101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11011010100101010000) && ({row_reg, col_reg}<20'b11011010101000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11011010101000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b11011010101000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==20'b11011010101000111000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11011010101000111001) && ({row_reg, col_reg}<20'b11011010101000111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11011010101000111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11011010101000111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11011010101000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11011010101000111111) && ({row_reg, col_reg}<20'b11011010101001100000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11011010101001100000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11011010101001100001) && ({row_reg, col_reg}<20'b11011010101001100101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11011010101001100101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11011010101001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11011010101001100111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11011010101001101000)) color_data = 12'b101110111011;

		if(({row_reg, col_reg}>=20'b11011010101001101001) && ({row_reg, col_reg}<20'b11011010110100011100)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11011010110100011100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==20'b11011010110100011101)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11011010110100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b11011010110100011111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11011010110100100000) && ({row_reg, col_reg}<20'b11011010110100100100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11011010110100100100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11011010110100100101) && ({row_reg, col_reg}<20'b11011010110101001001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11011010110101001001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11011010110101001010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b11011010110101001011) && ({row_reg, col_reg}<20'b11011010110101001101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11011010110101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11011010110101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11011010110101001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11011010110101010000) && ({row_reg, col_reg}<20'b11011010111000110110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11011010111000110110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b11011010111000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==20'b11011010111000111000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11011010111000111001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11011010111000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11011010111000111011) && ({row_reg, col_reg}<20'b11011010111000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11011010111000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11011010111000111111) && ({row_reg, col_reg}<20'b11011010111001100000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11011010111001100000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11011010111001100001) && ({row_reg, col_reg}<20'b11011010111001100100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b11011010111001100100) && ({row_reg, col_reg}<20'b11011010111001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11011010111001101000)) color_data = 12'b101110111011;

		if(({row_reg, col_reg}>=20'b11011010111001101001) && ({row_reg, col_reg}<20'b11011011000100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11011011000100011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b11011011000100011111) && ({row_reg, col_reg}<20'b11011011000100100001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11011011000100100001) && ({row_reg, col_reg}<20'b11011011000100100100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11011011000100100100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11011011000100100101) && ({row_reg, col_reg}<20'b11011011000101001001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11011011000101001001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11011011000101001010) && ({row_reg, col_reg}<20'b11011011000101001110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11011011000101001110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==20'b11011011000101001111)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b11011011000101010000) && ({row_reg, col_reg}<20'b11011011001000110111)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11011011001000110111)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b11011011001000111000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11011011001000111001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11011011001000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11011011001000111011) && ({row_reg, col_reg}<20'b11011011001000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11011011001000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11011011001000111111) && ({row_reg, col_reg}<20'b11011011001001100100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b11011011001001100100) && ({row_reg, col_reg}<20'b11011011001001100111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11011011001001100111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==20'b11011011001001101000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==20'b11011011001001101001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11011011001001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b11011011001001101011) && ({row_reg, col_reg}<20'b11011011010100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11011011010100011110)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==20'b11011011010100011111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=20'b11011011010100100000) && ({row_reg, col_reg}<20'b11011011010100100010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11011011010100100010) && ({row_reg, col_reg}<20'b11011011010100100100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11011011010100100100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11011011010100100101) && ({row_reg, col_reg}<20'b11011011010101001001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11011011010101001001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11011011010101001010) && ({row_reg, col_reg}<20'b11011011010101001110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11011011010101001110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==20'b11011011010101001111)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=20'b11011011010101010000) && ({row_reg, col_reg}<20'b11011011011000110111)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11011011011000110111)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b11011011011000111000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==20'b11011011011000111001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11011011011000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11011011011000111011) && ({row_reg, col_reg}<20'b11011011011001100100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11011011011001100100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11011011011001100101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11011011011001100110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11011011011001100111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==20'b11011011011001101000)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=20'b11011011011001101001) && ({row_reg, col_reg}<20'b11011011100100011101)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11011011100100011101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==20'b11011011100100011110)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==20'b11011011100100011111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11011011100100100000) && ({row_reg, col_reg}<20'b11011011100100100010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11011011100100100010) && ({row_reg, col_reg}<20'b11011011100100100100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11011011100100100100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11011011100100100101) && ({row_reg, col_reg}<20'b11011011100100100111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11011011100100100111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11011011100100101000) && ({row_reg, col_reg}<20'b11011011100101001001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11011011100101001001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11011011100101001010) && ({row_reg, col_reg}<20'b11011011100101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11011011100101001101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11011011100101001110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==20'b11011011100101001111)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=20'b11011011100101010000) && ({row_reg, col_reg}<20'b11011011101000110111)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11011011101000110111)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==20'b11011011101000111000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==20'b11011011101000111001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11011011101000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11011011101000111011) && ({row_reg, col_reg}<20'b11011011101000111111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11011011101000111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11011011101001000000) && ({row_reg, col_reg}<20'b11011011101001100100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11011011101001100100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11011011101001100101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11011011101001100110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11011011101001100111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==20'b11011011101001101000)) color_data = 12'b110111011101;

		if(({row_reg, col_reg}>=20'b11011011101001101001) && ({row_reg, col_reg}<20'b11011011110100011101)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11011011110100011101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==20'b11011011110100011110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b11011011110100011111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11011011110100100000) && ({row_reg, col_reg}<20'b11011011110100100010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11011011110100100010) && ({row_reg, col_reg}<20'b11011011110100100100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11011011110100100100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11011011110100100101) && ({row_reg, col_reg}<20'b11011011110100100111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11011011110100100111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11011011110100101000) && ({row_reg, col_reg}<20'b11011011110101001001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11011011110101001001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11011011110101001010) && ({row_reg, col_reg}<20'b11011011110101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11011011110101001101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11011011110101001110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==20'b11011011110101001111)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b11011011110101010000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11011011110101010001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=20'b11011011110101010010) && ({row_reg, col_reg}<20'b11011011111000110100)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11011011111000110100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=20'b11011011111000110101) && ({row_reg, col_reg}<20'b11011011111000110111)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11011011111000110111)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b11011011111000111000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==20'b11011011111000111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11011011111000111010) && ({row_reg, col_reg}<20'b11011011111000111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11011011111000111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11011011111000111101) && ({row_reg, col_reg}<20'b11011011111000111111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11011011111000111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11011011111001000000) && ({row_reg, col_reg}<20'b11011011111001100100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11011011111001100100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11011011111001100101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11011011111001100110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11011011111001100111)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b11011011111001101000)) color_data = 12'b110111011101;

		if(({row_reg, col_reg}>=20'b11011011111001101001) && ({row_reg, col_reg}<20'b11011100000100011000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11011100000100011000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=20'b11011100000100011001) && ({row_reg, col_reg}<20'b11011100000100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11011100000100011110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b11011100000100011111)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b11011100000100100000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11011100000100100001) && ({row_reg, col_reg}<20'b11011100000100100100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11011100000100100100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11011100000100100101) && ({row_reg, col_reg}<20'b11011100000100100111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11011100000100100111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11011100000100101000) && ({row_reg, col_reg}<20'b11011100000101001000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11011100000101001000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11011100000101001001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11011100000101001010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11011100000101001011) && ({row_reg, col_reg}<20'b11011100000101001110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11011100000101001110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11011100000101001111) && ({row_reg, col_reg}<20'b11011100001000110100)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11011100001000110100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=20'b11011100001000110101) && ({row_reg, col_reg}<20'b11011100001000111000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11011100001000111000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11011100001000111001) && ({row_reg, col_reg}<20'b11011100001000111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11011100001000111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11011100001000111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11011100001000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11011100001000111111) && ({row_reg, col_reg}<20'b11011100001001100000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11011100001001100000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11011100001001100001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b11011100001001100010) && ({row_reg, col_reg}<20'b11011100001001100101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11011100001001100101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11011100001001100110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11011100001001100111)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b11011100001001101000) && ({row_reg, col_reg}<20'b11011100001001101010)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11011100001001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b11011100001001101011) && ({row_reg, col_reg}<20'b11011100010100011111)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11011100010100011111)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=20'b11011100010100100000) && ({row_reg, col_reg}<20'b11011100010100100010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11011100010100100010) && ({row_reg, col_reg}<20'b11011100010100100101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11011100010100100101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11011100010100100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11011100010100100111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11011100010100101000) && ({row_reg, col_reg}<20'b11011100010101001010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11011100010101001010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11011100010101001011) && ({row_reg, col_reg}<20'b11011100010101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11011100010101001101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11011100010101001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b11011100010101001111) && ({row_reg, col_reg}<20'b11011100011000111000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11011100011000111000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b11011100011000111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11011100011000111010) && ({row_reg, col_reg}<20'b11011100011000111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11011100011000111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11011100011000111101) && ({row_reg, col_reg}<20'b11011100011001100000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b11011100011001100000) && ({row_reg, col_reg}<20'b11011100011001100011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11011100011001100011) && ({row_reg, col_reg}<20'b11011100011001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11011100011001100110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==20'b11011100011001100111)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=20'b11011100011001101000) && ({row_reg, col_reg}<20'b11011100011001101010)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11011100011001101010)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b11011100011001101011) && ({row_reg, col_reg}<20'b11011100100100011101)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11011100100100011101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==20'b11011100100100011110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11011100100100011111)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b11011100100100100000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=20'b11011100100100100001) && ({row_reg, col_reg}<20'b11011100100100100101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b11011100100100100101) && ({row_reg, col_reg}<20'b11011100100100100111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11011100100100100111) && ({row_reg, col_reg}<20'b11011100100101001000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11011100100101001000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11011100100101001001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b11011100100101001010) && ({row_reg, col_reg}<20'b11011100100101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11011100100101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11011100100101001101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11011100100101001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b11011100100101001111) && ({row_reg, col_reg}<20'b11011100101000111000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11011100101000111000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b11011100101000111001) && ({row_reg, col_reg}<20'b11011100101000111101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11011100101000111101) && ({row_reg, col_reg}<20'b11011100101000111111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11011100101000111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11011100101001000000) && ({row_reg, col_reg}<20'b11011100101001100001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11011100101001100001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11011100101001100010) && ({row_reg, col_reg}<20'b11011100101001100100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11011100101001100100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11011100101001100101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11011100101001100110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==20'b11011100101001100111)) color_data = 12'b110111011101;

		if(({row_reg, col_reg}>=20'b11011100101001101000) && ({row_reg, col_reg}<20'b11011100110100011111)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11011100110100011111)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b11011100110100100000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==20'b11011100110100100001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11011100110100100010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11011100110100100011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11011100110100100100) && ({row_reg, col_reg}<20'b11011100110101001000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11011100110101001000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11011100110101001001) && ({row_reg, col_reg}<20'b11011100110101001011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b11011100110101001011) && ({row_reg, col_reg}<20'b11011100110101001101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11011100110101001101)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==20'b11011100110101001110)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=20'b11011100110101001111) && ({row_reg, col_reg}<20'b11011100111000110111)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11011100111000110111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==20'b11011100111000111000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==20'b11011100111000111001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=20'b11011100111000111010) && ({row_reg, col_reg}<20'b11011100111000111101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11011100111000111101) && ({row_reg, col_reg}<20'b11011100111000111111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11011100111000111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11011100111001000000) && ({row_reg, col_reg}<20'b11011100111001100011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b11011100111001100011) && ({row_reg, col_reg}<20'b11011100111001100101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11011100111001100101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11011100111001100110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==20'b11011100111001100111)) color_data = 12'b110111011101;

		if(({row_reg, col_reg}>=20'b11011100111001101000) && ({row_reg, col_reg}<20'b11011101000100011111)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11011101000100011111)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b11011101000100100000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==20'b11011101000100100001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11011101000100100010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11011101000100100011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11011101000100100100) && ({row_reg, col_reg}<20'b11011101000101001000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11011101000101001000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11011101000101001001) && ({row_reg, col_reg}<20'b11011101000101001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11011101000101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11011101000101001101)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b11011101000101001110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=20'b11011101000101001111) && ({row_reg, col_reg}<20'b11011101001000111000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11011101001000111000)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b11011101001000111001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==20'b11011101001000111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11011101001000111011) && ({row_reg, col_reg}<20'b11011101001000111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11011101001000111101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11011101001000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11011101001000111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11011101001001000000) && ({row_reg, col_reg}<20'b11011101001001100000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11011101001001100000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11011101001001100001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b11011101001001100010) && ({row_reg, col_reg}<20'b11011101001001100100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11011101001001100100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11011101001001100101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11011101001001100110)) color_data = 12'b101110111011;

		if(({row_reg, col_reg}>=20'b11011101001001100111) && ({row_reg, col_reg}<20'b11011101010100100000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11011101010100100000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==20'b11011101010100100001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=20'b11011101010100100010) && ({row_reg, col_reg}<20'b11011101010100100101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11011101010100100101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11011101010100100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11011101010100100111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11011101010100101000) && ({row_reg, col_reg}<20'b11011101010101001001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11011101010101001001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11011101010101001010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11011101010101001011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11011101010101001100)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==20'b11011101010101001101)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=20'b11011101010101001110) && ({row_reg, col_reg}<20'b11011101011000111001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11011101011000111001)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b11011101011000111010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=20'b11011101011000111011) && ({row_reg, col_reg}<20'b11011101011000111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11011101011000111101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11011101011000111110) && ({row_reg, col_reg}<20'b11011101011001100000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11011101011001100000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11011101011001100001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11011101011001100010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11011101011001100011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11011101011001100100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11011101011001100101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==20'b11011101011001100110)) color_data = 12'b110111011101;

		if(({row_reg, col_reg}>=20'b11011101011001100111) && ({row_reg, col_reg}<20'b11011101100100100000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11011101100100100000)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b11011101100100100001)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b11011101100100100010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11011101100100100011) && ({row_reg, col_reg}<20'b11011101100100100101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11011101100100100101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11011101100100100110) && ({row_reg, col_reg}<20'b11011101100101001001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b11011101100101001001) && ({row_reg, col_reg}<20'b11011101100101001011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11011101100101001011)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==20'b11011101100101001100)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b11011101100101001101) && ({row_reg, col_reg}<20'b11011101101000111001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11011101101000111001)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b11011101101000111010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==20'b11011101101000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11011101101000111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11011101101000111101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11011101101000111110) && ({row_reg, col_reg}<20'b11011101101001100001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11011101101001100001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11011101101001100010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11011101101001100011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11011101101001100100)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==20'b11011101101001100101)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=20'b11011101101001100110) && ({row_reg, col_reg}<20'b11011101110100100001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11011101110100100001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==20'b11011101110100100010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==20'b11011101110100100011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11011101110100100100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11011101110100100101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11011101110100100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11011101110100100111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11011101110100101000) && ({row_reg, col_reg}<20'b11011101110101001000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11011101110101001000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11011101110101001001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11011101110101001010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11011101110101001011)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==20'b11011101110101001100)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=20'b11011101110101001101) && ({row_reg, col_reg}<20'b11011101111000110000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11011101111000110000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=20'b11011101111000110001) && ({row_reg, col_reg}<20'b11011101111000111010)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11011101111000111010)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==20'b11011101111000111011)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=20'b11011101111000111100) && ({row_reg, col_reg}<20'b11011101111000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11011101111000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11011101111000111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11011101111001000000) && ({row_reg, col_reg}<20'b11011101111001100001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11011101111001100001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11011101111001100010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11011101111001100011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11011101111001100100)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b11011101111001100101)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b11011101111001100110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=20'b11011101111001100111) && ({row_reg, col_reg}<20'b11011101111001101001)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b11011101111001101001) && ({row_reg, col_reg}<20'b11011110000100100010)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11011110000100100010)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==20'b11011110000100100011)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=20'b11011110000100100100) && ({row_reg, col_reg}<20'b11011110000100100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11011110000100100110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11011110000100100111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b11011110000100101000) && ({row_reg, col_reg}<20'b11011110000100101010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11011110000100101010) && ({row_reg, col_reg}<20'b11011110000100101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b11011110000100101100) && ({row_reg, col_reg}<20'b11011110000100101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11011110000100101110) && ({row_reg, col_reg}<20'b11011110000101000010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b11011110000101000010) && ({row_reg, col_reg}<20'b11011110000101000100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11011110000101000100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b11011110000101000101) && ({row_reg, col_reg}<20'b11011110000101000111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11011110000101000111) && ({row_reg, col_reg}<20'b11011110000101001001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11011110000101001001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11011110000101001010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==20'b11011110000101001011)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=20'b11011110000101001100) && ({row_reg, col_reg}<20'b11011110001000111000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=20'b11011110001000111000) && ({row_reg, col_reg}<20'b11011110001000111010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==20'b11011110001000111010)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11011110001000111011)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b11011110001000111100) && ({row_reg, col_reg}<20'b11011110001000111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11011110001000111111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11011110001001000000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11011110001001000001) && ({row_reg, col_reg}<20'b11011110001001000101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11011110001001000101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11011110001001000110) && ({row_reg, col_reg}<20'b11011110001001011011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b11011110001001011011) && ({row_reg, col_reg}<20'b11011110001001011101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11011110001001011101) && ({row_reg, col_reg}<20'b11011110001001100000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11011110001001100000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11011110001001100001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11011110001001100010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11011110001001100011)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==20'b11011110001001100100)) color_data = 12'b110111011101;

		if(({row_reg, col_reg}>=20'b11011110001001100101) && ({row_reg, col_reg}<20'b11011110010100100000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11011110010100100000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==20'b11011110010100100001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11011110010100100010)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b11011110010100100011)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b11011110010100100100)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==20'b11011110010100100101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11011110010100100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11011110010100100111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11011110010100101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b11011110010100101001) && ({row_reg, col_reg}<20'b11011110010100101011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11011110010100101011) && ({row_reg, col_reg}<20'b11011110010101000000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11011110010101000000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11011110010101000001) && ({row_reg, col_reg}<20'b11011110010101000011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11011110010101000011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11011110010101000100) && ({row_reg, col_reg}<20'b11011110010101000111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b11011110010101000111) && ({row_reg, col_reg}<20'b11011110010101001010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11011110010101001010)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b11011110010101001011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b11011110010101001100)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11011110010101001101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=20'b11011110010101001110) && ({row_reg, col_reg}<20'b11011110011000111011)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11011110011000111011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b11011110011000111100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==20'b11011110011000111101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11011110011000111110) && ({row_reg, col_reg}<20'b11011110011001000000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b11011110011001000000) && ({row_reg, col_reg}<20'b11011110011001000011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11011110011001000011) && ({row_reg, col_reg}<20'b11011110011001000110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b11011110011001000110) && ({row_reg, col_reg}<20'b11011110011001001000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11011110011001001000) && ({row_reg, col_reg}<20'b11011110011001011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b11011110011001011000) && ({row_reg, col_reg}<20'b11011110011001011010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11011110011001011010) && ({row_reg, col_reg}<20'b11011110011001011101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b11011110011001011101) && ({row_reg, col_reg}<20'b11011110011001011111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11011110011001011111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11011110011001100000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11011110011001100001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11011110011001100010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==20'b11011110011001100011)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b11011110011001100100) && ({row_reg, col_reg}<20'b11011110011001100110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11011110011001100110)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b11011110011001100111) && ({row_reg, col_reg}<20'b11011110100100100011)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11011110100100100011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b11011110100100100100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==20'b11011110100100100101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11011110100100100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11011110100100100111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11011110100100101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b11011110100100101001) && ({row_reg, col_reg}<20'b11011110100100110000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11011110100100110000) && ({row_reg, col_reg}<20'b11011110100101000010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b11011110100101000010) && ({row_reg, col_reg}<20'b11011110100101000110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11011110100101000110) && ({row_reg, col_reg}<20'b11011110100101001000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11011110100101001000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11011110100101001001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==20'b11011110100101001010)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=20'b11011110100101001011) && ({row_reg, col_reg}<20'b11011110100101001101)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11011110100101001101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=20'b11011110100101001110) && ({row_reg, col_reg}<20'b11011110101000111100)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11011110101000111100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==20'b11011110101000111101)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==20'b11011110101000111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11011110101000111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11011110101001000000) && ({row_reg, col_reg}<20'b11011110101001000011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b11011110101001000011) && ({row_reg, col_reg}<20'b11011110101001000110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11011110101001000110) && ({row_reg, col_reg}<20'b11011110101001011010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11011110101001011010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11011110101001011011) && ({row_reg, col_reg}<20'b11011110101001011101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11011110101001011101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11011110101001011110) && ({row_reg, col_reg}<20'b11011110101001100001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11011110101001100001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11011110101001100010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==20'b11011110101001100011)) color_data = 12'b110111011101;

		if(({row_reg, col_reg}>=20'b11011110101001100100) && ({row_reg, col_reg}<20'b11011110110100100010)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11011110110100100010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==20'b11011110110100100011)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11011110110100100100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==20'b11011110110100100101)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=20'b11011110110100100110) && ({row_reg, col_reg}<20'b11011110110100101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11011110110100101001) && ({row_reg, col_reg}<20'b11011110110101000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11011110110101000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11011110110101000010) && ({row_reg, col_reg}<20'b11011110110101000101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b11011110110101000101) && ({row_reg, col_reg}<20'b11011110110101001000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11011110110101001000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==20'b11011110110101001001)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b11011110110101001010)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11011110110101001011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=20'b11011110110101001100) && ({row_reg, col_reg}<20'b11011110111000111100)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11011110111000111100)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b11011110111000111101)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b11011110111000111110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=20'b11011110111000111111) && ({row_reg, col_reg}<20'b11011110111001000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11011110111001000001) && ({row_reg, col_reg}<20'b11011110111001011001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b11011110111001011001) && ({row_reg, col_reg}<20'b11011110111001011011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11011110111001011011) && ({row_reg, col_reg}<20'b11011110111001011110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b11011110111001011110) && ({row_reg, col_reg}<20'b11011110111001100001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11011110111001100001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==20'b11011110111001100010)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=20'b11011110111001100011) && ({row_reg, col_reg}<20'b11011111000100100010)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=20'b11011111000100100010) && ({row_reg, col_reg}<20'b11011111000100100100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==20'b11011111000100100100)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b11011111000100100101)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b11011111000100100110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==20'b11011111000100100111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11011111000100101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11011111000100101001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b11011111000100101010) && ({row_reg, col_reg}<20'b11011111000100101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11011111000100101100) && ({row_reg, col_reg}<20'b11011111000100101110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b11011111000100101110) && ({row_reg, col_reg}<20'b11011111000100110000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11011111000100110000) && ({row_reg, col_reg}<20'b11011111000101000000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11011111000101000000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11011111000101000001) && ({row_reg, col_reg}<20'b11011111000101000011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b11011111000101000011) && ({row_reg, col_reg}<20'b11011111000101000101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11011111000101000101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11011111000101000110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11011111000101000111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==20'b11011111000101001000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b11011111000101001001)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=20'b11011111000101001010) && ({row_reg, col_reg}<20'b11011111001000111101)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11011111001000111101)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b11011111001000111110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b11011111001000111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11011111001001000000) && ({row_reg, col_reg}<20'b11011111001001000010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b11011111001001000010) && ({row_reg, col_reg}<20'b11011111001001000101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11011111001001000101) && ({row_reg, col_reg}<20'b11011111001001000111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11011111001001000111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11011111001001001000) && ({row_reg, col_reg}<20'b11011111001001011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11011111001001011000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11011111001001011001) && ({row_reg, col_reg}<20'b11011111001001011011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b11011111001001011011) && ({row_reg, col_reg}<20'b11011111001001011101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11011111001001011101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b11011111001001011110) && ({row_reg, col_reg}<20'b11011111001001100000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11011111001001100000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==20'b11011111001001100001)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==20'b11011111001001100010)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=20'b11011111001001100011) && ({row_reg, col_reg}<20'b11011111001001100101)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11011111001001100101)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==20'b11011111001001100110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11011111001001100111)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b11011111001001101000) && ({row_reg, col_reg}<20'b11011111010100100101)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11011111010100100101)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b11011111010100100110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b11011111010100100111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==20'b11011111010100101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11011111010100101001) && ({row_reg, col_reg}<20'b11011111010100101011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11011111010100101011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11011111010100101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b11011111010100101101) && ({row_reg, col_reg}<20'b11011111010100110000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11011111010100110000) && ({row_reg, col_reg}<20'b11011111010101000100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b11011111010101000100) && ({row_reg, col_reg}<20'b11011111010101000110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11011111010101000110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==20'b11011111010101000111)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b11011111010101001000)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b11011111010101001001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=20'b11011111010101001010) && ({row_reg, col_reg}<20'b11011111010101001100)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11011111010101001100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=20'b11011111010101001101) && ({row_reg, col_reg}<20'b11011111011000111011)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11011111011000111011)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=20'b11011111011000111100) && ({row_reg, col_reg}<20'b11011111011000111110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11011111011000111110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b11011111011000111111)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b11011111011001000000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==20'b11011111011001000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11011111011001000010) && ({row_reg, col_reg}<20'b11011111011001000100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b11011111011001000100) && ({row_reg, col_reg}<20'b11011111011001000110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11011111011001000110) && ({row_reg, col_reg}<20'b11011111011001011010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b11011111011001011010) && ({row_reg, col_reg}<20'b11011111011001011100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11011111011001011100) && ({row_reg, col_reg}<20'b11011111011001011110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11011111011001011110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==20'b11011111011001011111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==20'b11011111011001100000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=20'b11011111011001100001) && ({row_reg, col_reg}<20'b11011111011001100101)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11011111011001100101)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b11011111011001100110) && ({row_reg, col_reg}<20'b11011111100100100000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=20'b11011111100100100000) && ({row_reg, col_reg}<20'b11011111100100100010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=20'b11011111100100100010) && ({row_reg, col_reg}<20'b11011111100100100100)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11011111100100100100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==20'b11011111100100100101)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11011111100100100110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b11011111100100100111)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==20'b11011111100100101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==20'b11011111100100101001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==20'b11011111100100101010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11011111100100101011) && ({row_reg, col_reg}<20'b11011111100100101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b11011111100100101101) && ({row_reg, col_reg}<20'b11011111100100101111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11011111100100101111) && ({row_reg, col_reg}<20'b11011111100101000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b11011111100101000001) && ({row_reg, col_reg}<20'b11011111100101000101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11011111100101000101)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b11011111100101000110)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=20'b11011111100101000111) && ({row_reg, col_reg}<20'b11011111101000111111)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11011111101000111111)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b11011111101001000000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==20'b11011111101001000001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==20'b11011111101001000010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11011111101001000011) && ({row_reg, col_reg}<20'b11011111101001000101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b11011111101001000101) && ({row_reg, col_reg}<20'b11011111101001001000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11011111101001001000) && ({row_reg, col_reg}<20'b11011111101001011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b11011111101001011000) && ({row_reg, col_reg}<20'b11011111101001011010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11011111101001011010) && ({row_reg, col_reg}<20'b11011111101001011100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11011111101001011100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11011111101001011101)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==20'b11011111101001011110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b11011111101001011111)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b11011111101001100000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=20'b11011111101001100001) && ({row_reg, col_reg}<20'b11011111101001100011)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b11011111101001100011) && ({row_reg, col_reg}<20'b11011111110100101000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11011111110100101000)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b11011111110100101001)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b11011111110100101010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=20'b11011111110100101011) && ({row_reg, col_reg}<20'b11011111110100101101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11011111110100101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11011111110100101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11011111110100101111) && ({row_reg, col_reg}<20'b11011111110101000010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11011111110101000010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11011111110101000011)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==20'b11011111110101000100)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b11011111110101000101)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=20'b11011111110101000110) && ({row_reg, col_reg}<20'b11011111110101001000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11011111110101001000)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}==20'b11011111110101001001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=20'b11011111110101001010) && ({row_reg, col_reg}<20'b11011111110101001100)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=20'b11011111110101001100) && ({row_reg, col_reg}<20'b11011111111000111001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11011111111000111001)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=20'b11011111111000111010) && ({row_reg, col_reg}<20'b11011111111001000001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11011111111001000001)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b11011111111001000010)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b11011111111001000011)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=20'b11011111111001000100) && ({row_reg, col_reg}<20'b11011111111001000110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11011111111001000110) && ({row_reg, col_reg}<20'b11011111111001011011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11011111111001011011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11011111111001011100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==20'b11011111111001011101)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==20'b11011111111001011110)) color_data = 12'b110111011101;

		if(({row_reg, col_reg}>=20'b11011111111001011111) && ({row_reg, col_reg}<20'b11100000000100101010)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11100000000100101010)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==20'b11100000000100101011)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==20'b11100000000100101100)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==20'b11100000000100101101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11100000000100101110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11100000000100101111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11100000000100110000) && ({row_reg, col_reg}<20'b11100000000100110010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b11100000000100110010) && ({row_reg, col_reg}<20'b11100000000100110101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11100000000100110101) && ({row_reg, col_reg}<20'b11100000000100110111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11100000000100110111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11100000000100111000) && ({row_reg, col_reg}<20'b11100000000100111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b11100000000100111010) && ({row_reg, col_reg}<20'b11100000000100111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11100000000100111100) && ({row_reg, col_reg}<20'b11100000000100111111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b11100000000100111111) && ({row_reg, col_reg}<20'b11100000000101000010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11100000000101000010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==20'b11100000000101000011)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=20'b11100000000101000100) && ({row_reg, col_reg}<20'b11100000001001000011)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11100000001001000011)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==20'b11100000001001000100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11100000001001000101) && ({row_reg, col_reg}<20'b11100000001001001000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11100000001001001000) && ({row_reg, col_reg}<20'b11100000001001001011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11100000001001001011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11100000001001001100) && ({row_reg, col_reg}<20'b11100000001001001110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11100000001001001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11100000001001001111) && ({row_reg, col_reg}<20'b11100000001001010110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b11100000001001010110) && ({row_reg, col_reg}<20'b11100000001001011011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11100000001001011011)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==20'b11100000001001011100)) color_data = 12'b110011001100;

		if(({row_reg, col_reg}>=20'b11100000001001011101) && ({row_reg, col_reg}<20'b11100000010100101011)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11100000010100101011)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b11100000010100101100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==20'b11100000010100101101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==20'b11100000010100101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11100000010100101111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11100000010100110000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11100000010100110001) && ({row_reg, col_reg}<20'b11100000010100111000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11100000010100111000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11100000010100111001) && ({row_reg, col_reg}<20'b11100000010100111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b11100000010100111101) && ({row_reg, col_reg}<20'b11100000010101000000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11100000010101000000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==20'b11100000010101000001)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b11100000010101000010)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=20'b11100000010101000011) && ({row_reg, col_reg}<20'b11100000011001000100)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11100000011001000100)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b11100000011001000101)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b11100000011001000110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=20'b11100000011001000111) && ({row_reg, col_reg}<20'b11100000011001001001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11100000011001001001) && ({row_reg, col_reg}<20'b11100000011001001110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11100000011001001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11100000011001001111) && ({row_reg, col_reg}<20'b11100000011001010011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==20'b11100000011001010011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11100000011001010100) && ({row_reg, col_reg}<20'b11100000011001010110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=20'b11100000011001010110) && ({row_reg, col_reg}<20'b11100000011001011000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11100000011001011000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==20'b11100000011001011001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==20'b11100000011001011010)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==20'b11100000011001011011)) color_data = 12'b110111011101;

		if(({row_reg, col_reg}>=20'b11100000011001011100) && ({row_reg, col_reg}<20'b11100000100100101101)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11100000100100101101)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=20'b11100000100100101110) && ({row_reg, col_reg}<20'b11100000100100110000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b11100000100100110000) && ({row_reg, col_reg}<20'b11100000100100110011)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11100000100100110011) && ({row_reg, col_reg}<20'b11100000100100110101)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=20'b11100000100100110101) && ({row_reg, col_reg}<20'b11100000100100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11100000100100111001) && ({row_reg, col_reg}<20'b11100000100100111011)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=20'b11100000100100111011) && ({row_reg, col_reg}<20'b11100000100100111101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11100000100100111101) && ({row_reg, col_reg}<20'b11100000100100111111)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b11100000100100111111)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=20'b11100000100101000000) && ({row_reg, col_reg}<20'b11100000100101000010)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=20'b11100000100101000010) && ({row_reg, col_reg}<20'b11100000101001000000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=20'b11100000101001000000) && ({row_reg, col_reg}<20'b11100000101001000010)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=20'b11100000101001000010) && ({row_reg, col_reg}<20'b11100000101001000110)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11100000101001000110)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}>=20'b11100000101001000111) && ({row_reg, col_reg}<20'b11100000101001001001)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=20'b11100000101001001001) && ({row_reg, col_reg}<20'b11100000101001001100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11100000101001001100) && ({row_reg, col_reg}<20'b11100000101001001110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=20'b11100000101001001110) && ({row_reg, col_reg}<20'b11100000101001010010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=20'b11100000101001010010) && ({row_reg, col_reg}<20'b11100000101001010100)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=20'b11100000101001010100) && ({row_reg, col_reg}<20'b11100000101001010110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=20'b11100000101001010110) && ({row_reg, col_reg}<20'b11100000101001011000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b11100000101001011000)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==20'b11100000101001011001)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=20'b11100000101001011010) && ({row_reg, col_reg}<20'b11100000101001011100)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11100000101001011100)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b11100000101001011101) && ({row_reg, col_reg}<20'b11100000110100110000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=20'b11100000110100110000) && ({row_reg, col_reg}<20'b11100000110100110010)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}==20'b11100000110100110010)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==20'b11100000110100110011)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b11100000110100110100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==20'b11100000110100110101)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=20'b11100000110100110110) && ({row_reg, col_reg}<20'b11100000110100111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11100000110100111001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==20'b11100000110100111010)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b11100000110100111011)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==20'b11100000110100111100)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=20'b11100000110100111101) && ({row_reg, col_reg}<20'b11100000110101000101)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}>=20'b11100000110101000101) && ({row_reg, col_reg}<20'b11100000110101000111)) color_data = 12'b111111111111;
		if(({row_reg, col_reg}>=20'b11100000110101000111) && ({row_reg, col_reg}<20'b11100000111001001001)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11100000111001001001)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=20'b11100000111001001010) && ({row_reg, col_reg}<20'b11100000111001001100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==20'b11100000111001001100)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b11100000111001001101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==20'b11100000111001001110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=20'b11100000111001001111) && ({row_reg, col_reg}<20'b11100000111001010001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==20'b11100000111001010001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==20'b11100000111001010010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==20'b11100000111001010011)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==20'b11100000111001010100)) color_data = 12'b110011001100;
		if(({row_reg, col_reg}==20'b11100000111001010101)) color_data = 12'b110111011101;
		if(({row_reg, col_reg}>=20'b11100000111001010110) && ({row_reg, col_reg}<20'b11100000111001011000)) color_data = 12'b111011101110;
		if(({row_reg, col_reg}==20'b11100000111001011000)) color_data = 12'b111111111111;

		if(({row_reg, col_reg}>=20'b11100000111001011001) && ({row_reg, col_reg}<=20'b11100000111110000011)) color_data = 12'b111011101110;
	end
endmodule